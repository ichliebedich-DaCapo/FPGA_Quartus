-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LFNw2v2agmn+JpWjEss5izyYmRD2i4iOhH5cPW6MuMBfCgtCXErC/q4bRnms99+WqLVfG2OnrTR4
a3dxSQqP0JCMiXmpGuzCSkzZGYowNqgUYrQPwWuT3Phcl+xBl9a4/VdAwI5Ri0Z6IY7RM4LHWLbW
lbWjmfFWt/FWT4WxaXCr27as4bQPbeaS1GBlBSldolu7Qfgs+U5kB9+n8AUTgGOszlcFFR8dJL6J
BkxWra4oO3O5Z9T/D3Az7A3UlAOEDFb7E6xr/7K9/vcRavp1wZuIqKFsWZ/fi78O3yGkKvaUa5mn
Mdu7z9HGnIm/kY+BOjr7F876nDa9yfo/9xvM3g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
nfHh9KyXzeZv8bxKMcyR0WkrLBUmemRx1ZMAZD5ci2DX6o7h9vac5bbCGFIfTikP4BXsl60vkqqK
HKagt2ulq62Tye0QCcqirt6TQeroKFhMBirB0tNNUljJb8G0KxHnAQn/JIuaH4u65Ggdg/oKxjU6
EhrLAuBlp7XemptfFQRM8b5mCn8mK/Zm0vyTgIKI7lZlEXwRRbnB8ZKwsN++dLbDl8EZS9vFX0tE
eU5tdCoL8rAI4IaD1KXM76tEOvb2jvFpF/nRWRLEW4ip2tkra5t+jNvHBXpt7km3EPpDHrsirkWs
iRngpNwuWkaI/SfBEZ5jCHk2q4zRIeNljnatzumtvi6k3WYybPYWmj7aHVOAUbg21N9TywZEQKVe
dFI9jMfsM2n8GbhduHiL6/eMbKoUxiIix15Es4LSjijS/BIDs+RYqgoc5xXpiIBotYMXnG6GODcm
GnyWSG1biL49/lRYa9o+uNBnwtD8ALojVj+/yBXOG78AaoDQt8teBZejoFkMqCCq22ar+fZTpq3Y
C8MouEpY1PHvWhOwzmarzeoqe2QLzM+Kgv2oQeqD7dExEvUxKvbEnpWipeaT9KHTJ+75uyM2FHeJ
7J6cNAX4Iurz1Y9Rlnpi+v2ow1QVqpWKUiXvIyA29CVsqQ+xBuDwKhceSwP+aYZ6lWH2eiz7c2Te
emkVjaludWqCj2InhRG3ytL3x3RN0RdjCs6DRrbuyqX4v9V8QYz8supKq/UNwLtUgVGKsizVxtY1
PUKtQmEULZgRM4N5WeNvzZUc/OTjFAsG42n3Chca7yxnySWyLndbtlZRwLqgsfmozTwz5iwRrUka
Jix5/YPuzzZizMvfIbL2cfvIEHa1tih9BQhM9Sq5JtWSfwPm7u+Y6aLXTF0FhftMQIVElqk86gCm
UlpWpnR8UVWH21gw4DcYb8drMy73GINLc8awYB2O49gFpWidTVgF2zlfBJAq/xPJ++igmxzKxOEs
85jwRDTifDhmrlO0EazrV4VO4h1ISGlRyTIpqpm4aV+w9a0Ef/RXz61XbiIcB2inGQFpd074EwIg
aw5h6zQlNbt4YOTJct4lzUcMEbhnrmK7UxItMYDOf3XKcbXRURZy0P+5V+G6ahJ7/ftp22bS3h2W
cQmr4sLA3j3b596VWtUuPVpNKwxYfiOuYMiyk47MF42XavQVK0eX8X1v8toYE/Mt0/RO8XElRROJ
SW7xjQD39aMi7ei8YG2gaP4rVi0SqNLJjqOW7PdzaEvJhz96lOKGUjoTYmRHg4lonk3UTHvoOSoL
6LoyaTMWWfXHME6nXD626OnGnxdcXoPfK/zyuceehoFniERkPU/ZXKXYZXuJmamsnAGLzLjQQfk+
LrkFtQwaGh5cy9rqCk4ynYkhpjGRtZynSZgiQDyaUOtrR2qfIDPG+YG0vd5DpJyQtSbUB1s1gP+T
7NN2eR13o/8qgxdiGwggn/ynPzN/x+Q4USLU/aS59BkEVDErA198AcqthFq611qvHiyjzxQSu+kH
G/oW4E0jRAaYfvz6h4RgE0ECZ+IJ30FyS2sqCuHwTU6BwlWPgtXMAjzVy/zx6kRaui23SB84xViy
J+Zz4CHl+uHBPhNnhnbSyy/O3GG2w0xiOwummK5B68XBLH1jpsHWEPYYV2NBj2FdeZ/wuEvIrnrM
ecTiQuwEe1ENg55HBPECnD3vCgauzz/8d0Lf6KXKCchEHHRjkhJ/1kCBmW6VPzFBgNjFD260KQml
DEypxwhDUSsiZZOpSaQ5Gg8QksaoKwJi3cxINr6idVSvXeASgW9+xE2NC+bUfAkowNCu+OFYshoH
hIBpKWnt/mmKJmGp4H3mBeJm/F29EYr0oPZPTENV9GfTHi3EDIPbk+/lg6wGz2vbbhknoe1bbA/t
/cqw6Lb6Aug6gUs7W/9eNOfx7bT+OhfcLiF0wNcGRXSZ/HA39WABvdKxn/izdt+ab7DMg5u6r0nu
EBQfqhj0h86YG4XZPhKdSdUF/5pQfT80zA3Mj+clrq7WSkquufc9jhiBmAFmMFQvBXToBfKSr6P6
eS3vejnqYcs2xuZsByKyJmh+grzoJjboiNemah+Zq9BbGby3pCfDD0yBup0ZgS8elgAhpbkGRPQW
aBSgrMAZk1VG7GgA+jYsTvAZvktA20B8nWd0urOrOM5x7s9FSMP95s56nUKEN9Nvm58ndzDzH+mX
hlItElke75uV08YjcmHktzE+RHlPZNIOegkNE7iVH4pMADol/kwwQJTFObBe9guSuTQNi6au2Q0+
sThwzTa0Dk6B8jakJXnCe6FsZpaQMqi4mYDjw2EJyV93pJUakNWJ+4mjFnJy3bAoQv07U+WhVtt0
GnI47eGF+sdRxei3SdJCSmVd0hgPBIzuwl60RuckcFWHxzromyyao3F2gsIdQKciqncsOVWoCmjZ
g4mjJxE3Pz0l5CZnodX3DzZ4SiOh26BiHg8KYHyy+MilIlP3f/LWZ0cIRo1U8guHWkv4w2DkXJe2
MLEDwaH1QMrAVXmWzdXaWr7lBZ8JWdqL1kCkHM6/dpGP3mlnHCmM3X6YZldZa1GksQS5F/eYVsEM
uwos+emKbt2Nps8n6g5D2SOVmG9S5EKv3zfBfNKRiWtECfvPWJqykTsx4yrXKvQG5ovtB17jicMA
UeaFAFfyZxJx9NmiVEXJjMkuRyRqjbmWF3k0u3wIfas2M0J35mEOji/4H4Ser+OygDxDT1WfAroE
46vdhjLi25Opjrc5zR6GaGyoVg3tY//Ih2aqBP3Q3BWUkWbsioJMclMok4HQZeTcyRGuXHZxf2vj
kIpiBOK1OJoGP1LM+PXbrXOLhDHjXknyUxiBuWf2h4htB6rsADSmyVziSiT+syi/3UYdlWjffkQy
4+Ofh7GySH6x5Z2p4nsGLXVXkwVvpMR3cerF2TdiG7Cq5FuFQyRgq8XFdbx1Y5MlGcKm8nQ5QsRJ
8NAeETihd82hV1yXo2Eb8YPwXuLVZ+CzKFC7UFJnDxm+2kZUa2EexGQ88JqlNxRY/D52ABHwSy/W
qed0UY3cx/rxlzRvW8yTQyc0VJRTlvnNxcvAyeR8RKBaITu7057obNgExvVTCPHlz/2WJ7Sn2wZE
zerDnSb8xLmAmRh1ndJFRxx51YR9oZkLjAyuaMfRqzy4C/ZUeiVbzut1cK0uXXmYZEDZicfnZLw/
+Ybe4aXEGeU14MEZtlP9aZTmmXOZmhVi0xLlM5V8ZIqgfWj/VWvLfw+6WLTiedlw4OSlv8aEvUgI
/Le9rfYuGQP3y3FzUfGNC9VoQEsCT5cPUVMS52YAyn8AioO28OWm+CHKp9s3wI2d57SsshIMouDV
fscKr6Au0O0j+UvaqMykCe1Fo+0KDQE4fPEs1n5fSSBYivTFge9aBOZmS++ih+mVe0QkIasr5giP
3Ne+Hrb2j6/IrZ3kHzgZWDMaJPe0/b/RNXK7p4G5oNecd3Jnj3jErzUwxC0FyTZVI14M2reLactb
DfP7J+rEJAZTlgOmQM00SlxhOHglxvyziUc2Zp0PSDHkOZ/AiFcVdH6HkUfwxtocCxpvjU75+oZU
VCddTqUOS+Z8tWYQvY+QLiurnEZLRIgp5iIKNI77zbWlx4M/kU5ChVtz+we7mj6UmPTHOZ/VH/bt
/LajB1qBbFQYCikIlMyoLFBA+t344IXGp3ouGKcM6n37TvOkagbJB03Rqx3mUcxQIkghlu2jHrAU
BK9ZQZvSeaFvYo08pGckqKsbO90qArHryvH56qad/SpQKYShSW6Z5ymKn/KSJ5z2rOLUJsy+aGgt
5y6/RLPUB8zNPyCuUxfRsRTgShj4h0l55mNsUoAyecgXWM5HN6R5TNewxdCHWXburBeIrNncNoL1
RxXzYWaCq0UrW3us62xuKjtOhGzPKzNtxI8RHCfcr/dArZI7KIMNg7p86mNiJKoc48ROWX1rInHX
8F2/ZcD7HCBaWXNgnejRujC0NxUJPdoyTRyojqkxub/8R2NZxUMgm0Q47ZulvS3vvxBJ4R/j9DdX
q5ND6Rw7tJlu9CAKpA1tFBeHarY0Ecw2MlZXJSnMV29Q7DNiu9hmZEpulntf3l0zqy7ncveuGXTJ
QNOaWuP7usP7dnj0mH2pnV8WGdH9nr2enEnFL+pm2xaJFDZfr2z+CRfphladXwG/pnu0W8j7tqFp
XTPISb3MdbVs2GCV2QajG+4HUzkBHdpI1rGMWya+ZLYqw8OIWHvKoM3180x96RXV9ROVorxGd4BX
3+N7ujZNjMJylKLflZhNWJwmR96MyuISGRChIGGsc6Wa+kIlMMISBtHWHSSZKnsEMoGXJ5Wu6Yrj
uS/famo7tG3nQbOWBgv3cCnRGvh4vIN7jzcs7RI32cMMi5N3Sz0rsgmD80sw0JMudkHih/3v+RH/
nrIa8it+NzeCWhxngbhkCnzlf79DUPsJJaKI2GohqGiC2+BSVwV5MOJ778nFJkYSlT6XkDCe8njf
oXNSWqDdLJon924S8F6w0/ZyjYnEUFm84d3CxJvpqGF27SQSh4pYd9Qrojh7WsQ7RPvmri/8EetM
Y1UZtgazbiB2ajat8Wpq3yN/e4X5b7aoVPrw3H1ruCT/ug0a67RDpGQavO/ymdNQMmJXieS2zoUy
QqvK+irFB1+8vm74eaCBYjnrNcoBYKoMWWF5WsaXmeP3q0wk+x9tMDO04T3x9cgzy8ezvRJnq5Ph
ZIuFpeeq2G2dOj6uwE7OwrzsaSzmPZUos2khn1i7O5COj017XDhBlNbyeeiwtzvVRaiJhY70GC76
eOhT3CvbnZzZetaSPe4L5pbaoOfeWnMO9Lph3FmAtnhdzYw+QKs966OrQgk5RERIsIV0MMajWyNV
bMOZNU5zPLqpZzp7snXfRyR75z9cRNVMcEx4eXmSq50UwywZfPpbVt+d7t+POzjqmaEli4ukxAWM
UBbkp4fR7Wlof/0HKjQ46qvu9gds7cUI7yDhvP1J0WOGbQyISO7mmbA94geYz1XjeK6mELJhzyDg
SwuX10KGKtwZ8ocpNPhs47mJyy5UnHFk5Il8UBAH3gSncbK6WYOX91PsWcZFwFxkFUAcoRPIeH+R
ahOsJ3hpbeMav7eIEVzR4R/CAFXXq6D7sf6ouF2bwTzlBOgd0yaBXe9DDz4mGYJfCHopKTLY/W3E
9bLZ3kFGhqKPmDMydS+cYJ1xuPBi3A/6voySdKREwIkO8M5fFc+fXuBs24sVcbZIG3nFMhqM6d/p
e5gk6otnqGr7NNoiUxMZ/UH+y8mnzuGWPR7Zwq9hB7PEV3cWFm8GtsfmBOBadsNO309lto+bw7sm
9LcU9UNBmmf1KthnB4kACK+q4qbH5CTd/nhvCjfehG/NNnVjk5dyxqVGLZEz7OJxDfduWlmByZsb
qP7CAO6WG4wY3fdNDEm0p7kmnUAGCmbQBbQ33hfF0+mvkrLa7oA9XnfSTflD05whNCYtyl76v7da
8IblIGH/uGm/OfrYm8K6HkQHs02+9f2KUKxeo//Zv9kOTwRUi9cnqR2SGr+8AO2BnVbvPXmLRJtU
Qps3WG/O19k6MmLkxlASBN70CX9Qe8naLJxbhzVlv0Pf1jPo94wn76gblOech+Ma+y/ChKCD9jTW
tQ2DXccA6qkAQxF0HFoMX0/BHENZWMpVoaJpVXQOLaIcTAmNZAE63O2LXw17ukLO8oJaO169at2Z
BVOUJ224TltgPrnynA==
`protect end_protected
