-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I7e7c/3YgnVpnGB3+pfag6trbXN6989WHVGtXnWZYSZIZRFnlViHij/PcO8fPlIq1qEDNpa7INZH
wmD0jLBfYPfgHYGdWtYDG+28UIaNXRczG5yLRLXi8g9sRepfdI4Yi5kB5aS+7VHiKRBjcp/oWkFV
IJ2V+BVAibosVfh1ZMa2dYDxNrkfix2oZKsyZKZjMOrOT26A4uU91riiBd4BtaMZEpThY3Eoe74j
b63J37DN/stn8K8H3zAAdoKk/f/AOz9/MJzehfYNRedtxiIIXmAZEZZNhkFgXKh3qyQeiN2icz3L
2z058yv2j8XKKLxgTOfDs9l9ax02b+osJ/diWA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13920)
`protect data_block
KbT3QR5ScxbOr3ZPwZ7v3VLDWV74YL3zWc9JGaHWe3dC/Kqw4i/WmPRJOqyxD83atuu2ByPTGO8v
IF4mbkZX/ZRoSX5B1HYCRnB3CMo/OVaxAptUzDBA5x4RtgfdeYUAd1vo5FJaDKYu3922Fdr2CNXc
vJk8g3uhllD5tPa6bPFU5bGhcNXxevyxXGIAJFWT/M4bec/UNuiCrOgGnm3jY9p6ArcFhM8wW4s5
dysZ0gBSt2fYjFN5YP7hv2BsZbgP98ppJtbV0AFBSfWui2LKUtTWpAM+rc0tsfcnQHarQ7r1DPT4
H7WIqLcR9jWkVHuj3vJblTF42LpdBBO19KHYJFGfxA0NJy5QlACjhhG1vLIJ3ZYGm7Fn/jYHYlkV
WV3niLwZrIekOqNdNFZrOk6frz+aSAme57ndcCCVKpfS6dXBQycrJ1Jbk7300GDkzkY0fdMEl/Az
RR3mG9h8z7k4Kog/4fy/QPK5jSqcTNkoXJKqOa13h0v+e3OFTZtOzlp91zGKUxO9xIRYi4ypeSaa
y0mVhiojJN9GIqxn9dZ/Z26c5d4Wqs4+WDLPuNaJCqqKpBqtKzgFq20MW0aFhFpEobk09rY1NGJQ
+Xy7BeAN9MSXGvAVYxeti7n/5GHRqwh6VRotLsjVLWpbmDuJn/GRt7M964FQUDWam8tDXVooJODm
8/2qccRWae0eXfDnwiUhhDDWy5W6ANjricmw2w2YTf7pbt1GEIeXLD/PtVmydhmWl9UWmrm1A+B+
ahIqVAQ7RWMxVCSrO2khXCLfJYJi90OJ9rKWVXeIwX7KOHI/4ZKwPIb2KKUJ/WfVVCp5tP/YuVlV
uy+SJa/uv/8EIhfIC7GDjeVY4j7H7bgtmzd+b0lqjzrBK5vdyXDPrgwzSsrLL2cfadK/utEsyzQk
hZ9gxQ+q9/Uyhn8JC2aEVv72HKdUG6Qp+qxozB9d6KkomkNHjFn4h7079dUQ6S0wJksgueR04zNJ
oExxIfkpr9kByzqg+oKO6j0W0oaN61HVOgLDEsPM8INrlqlaKsA6KB80VHOQH2G+01nTXvpxAWeK
xIKJtSfsoo9UpR//VWDDgRWEfP+JNERCDZSv7Hffzi9glpfFOPqbg+BL3Wk/4g8J8hzOZYSXo8kA
lFf6stYzsziJC7cICZBSqusQeGqkf/JYBV74jLc9klCzvTp8GwtVZDiUOC6cLkNmkmVSkCQKRUp7
xjg7y46+gKu7KmbyqGoIy07/J9I8/PC0A1LjJD2vmwhZPLjYd2LJsIYSH4/fGZetYolqpLMnrzT8
eCrCiGHn1JCu00a8u6N7xr++izYa0+ComOW/8BoNYoZOUFX7YCOwpkCyE5dSaF/1GzViIlQ/jyPu
Zj1l9GgiOE4CqkvGwG+GFubZ2Z5gJhEvVFgwk8GqdjZD9rIiddpqN/l26ukqaoqyIDKpnvXAzJnY
2kJkbuWl8zawXA7ygb48NZui1b1y41PbnQoKBGO6xYQvyvJs+h9FFz98v4hsB5K9dnqCl5aZfDSC
yukvcygQ9vbEUY8B1l160cGCq+aMwC8FpIzPOdz5djYypcitBeei9x8ucjYr+KlxbRvo1GG3matd
hWHMY9mmkWuT5Umom/dl2RI4w5KDiU176I/uTZAZtPNm21JUQJCr1jheN75w2O802BgnC36V7alh
id6GVPbaDIwlUoZggbG4SvGdOnCJy13RNiwARa/SLyhmYbDCBLZjIJLq913//xQZx2XghZ0oCs0M
aTTXXtYPNZnfjmLOqp0XjERp7GrvUISxgUWATHDQ1gAgttlYSwBND/gJLRm6PO9MpC75eIxA48oD
M+pfTxRVZGVJ4pcrgWsukshuZz6tw/TK6f7aDrzokN9xbbzfwqDD6TX/aUWr3P6PX637TjDfzdY6
TMIZ9xCurFeU0pzHJhVDRZ1EtVPwTYjO/Jy1WrBumucMFnwPrtRPfA11NwVPWjQ/GWCzCNPEcIyo
qBDtZr4xW4FMLyLk4doAK0+2Ag5KMta/V/yVYZ6KWeO3fjUiJ5Z6kUv5pV6QKrqpFbGplu76ZUUz
7xE4WFQe5R39Y3LEOSmvmHhW2qu88oh8fsknFJYVPqculfhJjbUreU1PZmbFZO0ahbwaYC6GSg5x
FJ4srp5tVw3SUXv0vqsESIz7MD8O/9Qeb0ORi3nwO/HPVCMEjKxNBRw5P+zG7R7NlH1mjnxalsbb
2C+UVRak/I9Zv9aEDuhpIZa9xq213/R5xp8htP1OGZuTFR9LZwOFptAdOyd+zlMV5lsLZNuH9X8j
iuDT6z834vvWoZ+AY6j721Z3i3AO8kj8nu0vBnq+rZ09A5LrkIwPrXZ7J+mR2FIP58XjTJwyhV51
e/vv/v7QKmpjdX7NZI9YSv9UhMy1UdXr8W9QodYxEs90+or6AtGp6/vlXz9nirfno5zNHEbrh/lz
Wf8S6u9MCZ2YG8IF296ReYJlyd3U9edfy3s6iVFF7XMnWtm7ee2ARRtaOVwaUVn1QaiZ8v/oTUoF
uyFsIZltIWdpF2ASGmCBs6msWTfI65W5WIO4O6xwAMlchOY1mMaU8jNj0xTn+EUXyiWHKgXhyLWt
cAuM2bDRvBwbJir0PfF5z63NN7Dxyni9fkl84TK4P27ExG3ClWpmQ//YK0kv5uRpw39x2FoSBlLA
qh+sbmNV+AmZiaYcnxBgWmHpoj5pWd/GRkmoj5c90U/dIwNAKwymeyLi3YG7sqCl0+y+PV+qzS8c
bKNJEZiGCmuomM5TFvkBq916ycxK/v576vUghzYd01e5LJvD6yctLGVcA/WpAmLP8hjHy2hWR3Xz
MzEAyBnEfo48dtBs8ibGHJ7P/RpjotOgBvsP4xKl+vGuNgRJC+VBC56UgpVOfa6lbxdExMQwl8pn
y70uRkrkHOsh5LUhenVtoAIReMJy/cUBmpKyzUvQw+1GEc0WDhrT7HWXfZvitA5S0GVJv0mloG5t
wea4DILgB83A4qAJZWTQNWnh2tWzzbePpUL6qkY9xUTXJteJVOZ3zZw1ozEj4Zk0yqeIP2V0uhk8
WO4PjIotbg6Gh/k5oGD+22p2VKpG99O76LECiSE/Abt++FezdDLJhugqZqL090VkOALDarT2eOCC
BYdIBtYCcKTw5/gajAHoy0NYorkawFj1qvxx/hvii1D6CHKk/Kb3wE9lKBKilwzF2ngZcHaCwGWL
TWFKpC6WgJUiUfxJOqwlymA0fKtBRwcLINkuamZI2p2MQaxvswOYhFISnxqj2qFprb31BExuOind
Gy8m7lKBcFcPGMwt10YlDN9ZIJflL+H/gHlpwzJ/ch//Ply4dfs5WmYr8FYFUQFNq/iigBhwOfNr
WjNhl9IYzyTUGadBoxL6bCdSW9apyhjZBC6u6b+XPAyDedkrG4UetM6k4qwG0gvp63uSXNKnKt3u
U/3hetLTF/QvAYxb3YpM/uZIXgJZOlyEO6bgjNkZaSiW36kzlfWBHs2p8pZr9ojscWegajMla0tz
G5fRcs1SsP2uHKpUbL6NBV7IlyEEW5It2le5x1AmwW7KIBZiMJNXXQLFtl1VVJ/c1prOdIXl9GiX
WVFbWuVgxD9ToKlW467cB3XhDUqzbvBBzUNx4JWN2gEf7p/gKMMip66XGNxPdZ5bk6pRlV4Kin8P
UeikzYcjzuXfGe+xLhYqjMDzAvL3OUC9ox7L4vnFlFyuhasZoxDGCerTA7ucKnjcxrHmSrrMzeNj
NbNlCZ7PWB4v+og1J9cmijaC3oObk2EwkdjWmn0OrcF+8RdtqPIhTRiIjwYKpI+0iqtqT8OTMCMr
00Kibv49d8+CNKJXVsxWhfgWJci1hkRfipzJZP029Fy1nx9VfeJeoVF4E0GvH3pwsAIkv0opOTwA
L5W7an9NzBPgm6OC7MkdxtrW/kSQOlYiqQR2jhC6Isi94Eg6GvLOuyYmuIApk26xKbUC5rUmFuGt
bkNmlsEvjXBPVfoRXUdXMrh8xG1K1KoS9O4GBAHv40zpHSeQDPzug9A5nkClZhqenO1NCAZX4JSV
KnqUQ7z2cG5PPa6cvcczHidB8H0SGPvfwdw/cZ4kcxDtDVxm87PrcVg5uXqPO7SJ0ggSmsPnMEZK
EnXryszUe1GBiZRwZ7QuNsgp8s3rz+1CyfaNQVktn8/1+7ThNKkG/WU1LVeLR59/1I7dsDWSM83E
23YW1+7Ec+29Ufw7tRZBTlBmkI1b8lEzuqsZbBohQV5mLQrx9mti4jZsMVmEXc6TYnPL5i2yyzfP
edvWLuwOXLtt4GAmdbz+rrq8cenrI0VjQ2kPA4ygfrUTIPK5yp67kKf/FPa2NZvvni9olPrtCx0j
F0IVA6ImpoOuVFWl7J6Dy9jFHqB5bapat2UKuCCJg+cZdu+ROqVITHV76vgtqRdWmDVjQxfL48eh
cX51vSLioTYZhW43d5B32TgZi4hBw5sc0lJmlcf1FJGRez75DRgXHeOpyKxFXM7qU+VAiY69m8TW
PeeuvGBYQoEDyf3NkYxnfc8BCeawayPSOPVjQK8Yb4DvlYTEVz/35OKxMY1ObYUh4o7c4iUD1wiJ
j1Q0mQAVpcmDpuFgeTGqbKgvPuE9LndiJVbVlcfPb4zHOiXnCouYCkfwjLNXX2e6uUT+qX1DeJL1
UeTvoMmIUHucH0YQv57TanLwd1ojvg16xAhdn7dacgKzQPokgIHGjG8yFPkRg2Y4nNjXsBqn3cmS
SxXivkZzwYb0fWptW2gA2Inso1lfowPWBzzCxk+TEtQwxO/4lf1UUZb++e6Z8/UYN5MGrqX6HnrM
eMw9Ok5C3gFtMzdu1REqotxbj5sqKKygBAV1+2IuuDWQnQ96EGFeeQvU/F9nzvIJ/FCY8zwot+BP
Wac7i6lASnLB2mMW5k3A6SD2DEOJ9BXTki6DWcgwULo+LbdUOu5hXIg4uPJ3SdxAvpBn0/bq/qZ3
T0XzIBIXc8IrP5pHH+OC/K8n+pXJZ/XFUiuc1TNVjqoDfEMTyHPzEQX2l3cKkE9TUiFUGb0mzfwH
D0iprkYIftJfZdT1hnHlH1/yaK8jBnL0OHptOd0WmikqTm7AlQOQk0HiIXUvN6Z6VBILEOzT4nk6
k1BknQIAKNcEecWMUr3p8nq7HpRdyPMbOr6fzH5CGdHw0ShWfWAFyJIFyeX+BtaKR2V4kz8ihfZP
q17DDOH8WGBq6/BbuLaSZx+By/rsbYr6fhyLI/da2jJqRi95jzlEZu3+ffNySROjEbQNQfZWQjAN
LR/PNlipp/AvgwK82BbbA1VtLb4Z8qYzECd5lIBhMHxf/m0cQ3i2dgHa+d7fLfaC6XTNbac+cb4T
LCTzkqPSR2xK/cLn3MdHCX5C6Ank4RWhGSPaPF0/sHk55B8Ylo7iguouj6rm9s7oPVRdiAWyRHwP
m+JEh4qLhEdjX7SO+5ymGSPnWAdSexTZfgJ9QWYpXLBDOpOAlaMO3N8w7tSmKQmML44JncXsAhqu
hxtGmYTKy7xNDEFqhHjC6aivmhQ5yi1QB9Wt3Qe5O7H0sNk9KSqv/WOgsgHz164Mh0FVHYbC+0p5
LKhzx7+lTK1nD2augL9/0pl6m1AX/WrByRiaK3JSqjJ0oOJIpkKJdyPjn+iTCyhAI9MWhjGkB/30
sOFyjWunRBvV7SZbNGI7+NU7N/NgTnLi+RfoCdk7oflA3V6YQHKAHiplflEATNIfavoo62/ss7vJ
cYFLInAh0Vb30BmuGgX21Sfa0mWJi+qFwUpPgEPQhklP9YaRyVhfCVFD6O2iHfUoHaj+uTEm2K3v
VFCQBKzFcB3igNcEIaCFS4gXKmCXkOwyM3Wyy5JWCMQr9EJCpdz6Sm4CAG/SbCxBaHCV4SX5gdz/
uh97HNh4EYYJUknYSiSpAnlrtkJMiTsWDNmJTNNFqQNLw0bS/iANRYKtWhoEHjE+hatfJBPuaxfK
MchZdvmTgjYnyhBBdZ5nkg/+1UmvG60lSGNsfyRfVGoI6F492n9GAQdLATMJVnBKyOpfqcVX24K9
+eQ/3BrA9g+UxOgI3EBX1GCsg3KJRTin9ArWeAtasCQK1H3MoKUuEOZ+KDqMCvdpEJeIPsVgp17R
Ho506XX3jWyEd4+hC2Q/GkbQqdsZXlZRbZo0nsEF/cqcyi7nPLjScwORfMYDU6VNGD+mW8KQZP6D
ru98flk15UHQEekyBCHk6XcX6txQX6mHBdxUNyqiXJxHqNSN9tvwugi356Lu/L0q6ODbZU3Ev+Pc
IbaCVZhyjT1ZZgsYG99LwcJSpWUpPioLqM1oiouBu8GOLCt+GA+wfBv3AAp7fUnsZUg6AnVQDh5E
7g30QIKdosuZDPgs+IThiUZtYiG9ZRcDNhVubzfEK/5I58hA8NsjPAjKdMNBPLpPX0GcndhTHMoy
F1DmT6BfIAxwq9aJzC345hV15lotVyXOQiDlUZLuvbWDYO8hJfs9MXOmtDrypUJx2SjPpojR780I
/ABqRJCb6D/BXdmMcMaSnQJqe86xGBlVMk6ILNny8bBK/CIyUC/HpgIkQaUyHQSDRRPSMlgcdfm9
qf9tBQx1cxEjjwBy9lyluoTuHf6EfzteG3AO/RR1NNyCTTifL6MvfNBBq+0SOsiKDKu8m/tC+thn
YRJKMM4ewWbXyZdXCEKFKh4YP9MgGTAaly4dEuKRWl1ydkc7frO9LXQ6P7+wMilzqj9tyu/h1ZKv
F2bjUC6/O6rtVgJbjmWBOVX1TrclNm5gIGPwyLjbJ4D+ZobLKOiGh4n1ukGwxBFbNPNi70rnYTcC
aGGWPqgN/5xEycMMy7TsGDrgGye5DGy/vzYaMKPrjTxgynMBeg1t0YXzsVFZDz/mem7EjKrBbb9X
qjeKQw1kvtK6n009mvGJHcJgYS9VVAyf3PtiIt/Ai0UtC6EoMBcvPtzwFXONTtm772F2nZhOYvmQ
9JEm/xalD152p6JXi2tU5aOYepnD5Y2yoKXXecDSh1LDvVhg1yVi1Rsaw4ZBg9ngTUN6JfP/Y4aE
hGbjdoUQ/9EmYUBgqDw7KrDs1Tt4bMH3tRLP05wMW6jPUCmwtxqHvLHrrY09qui90lr9jiaBa2Lc
Y2Z+fx38ek4fG5Fh9h9xLeDKk3AFcLBi3F+UACV+WVz1aGvf3Es93w0QxhiSl8o87q0TH4UPjtUl
ZLaW+fhfermQH6FDX6I09nB/PfQpMZqs8fNR9ijtogwfbvK37e+acv0ru9XO00r1VHs7oD7zQ1xl
d/Ll2Blmw/szJaMGoHR/Mt2WtYyO3rFHAZji1aVXjzpT2QzZOR9iJrb3RTRkEBlA5cAcGA/sZGNx
GyVr8A57FGLTEiFBadfpYXW57nprs5Z5CCc0Z4VkYVsBHOaFfg4PshvAgToGbM4pv3r91d8j322e
g2obpLQnYij+lk2G9zEEric5xZLI+kwBzwOy8BmC59ktGsnGjg6viTXIZDzgy2O9WVHQ1cLiGLGr
+wXkt/awHf98gXZJhbectvvx4m7/5HQoAbZt0K57ptNibupObeuaiap8qfcypd5WdNS5UpmG68RA
Pe+MEqsvfoE5IUK3vzOnOWg96F+H4DTo+RKucKnJaNc7DqBIhfKMQD+8nLoTvUtqiReFgrUL9LIh
lKQUrIW4+4u7HTFo8xU8MPYFThGfSJg5o8Q8Vd7B6ucdykb1Cr67M/Q8+W7wVc5UMIn+adlri6wD
EX+fxmv/JcOhMk+n6fhwfoZSuF9xx919PbnNIXgBoijVhN5l8j7A/AqdX8WWBO26F5aQoneaGBMv
WTzPc6Xx3Kanhf3MUrqluXdHZReVSxMhy25Ik9mPvEdh3HxQhTu6Th01o6UHBVXYVLGFJP/xqAFP
79F8OLOEFl6uXgWGnrfG8D/cresHy4rlfAvu7iOHY6DOFTiqqdHpz9qRPHGZzFqTig+TMIyBCxBk
SUHBI030SN7bLOuSJK9/X76XP/qe3AiHoYH5Ihkm+zesdpBV9/SIfRzkLpJi2D3jIqmf8r34Xv4X
C9khrO5Q5BaWJ1k9uWzGT/O8QOTGDk7E0/CyAt37ysFCwDVPd+l+DCneQ4K3y/yVxKfb51DPfAig
cx0BSCXf2VcvTkH9rqp4b1Qzzdwi4aD0hXI0yY3e3Eh6Xnlgy/GRuMY2EnB6b3GdsRLtHBFDKbHk
+YhPVcxDfTVA+8XvOFgaZ3Pf68bJOhaIpZ241Ti66Z6XFkT9yRd77xRxW/tAoYYk/fSETmf+c2o5
Zer+sTgsOThronLbFK8VIflQzz44XBq73k0Qm4L7jzbo4KmPYPzI0lLrdaFq6IJu0VbF9hN+a2/k
JYvkqho6MwiiCyuIK7K+DW7Nvub+nceJz4YachQrWISXT0QfbT/nuAMLNgtIfOGva6bPOvqpX++m
YD4dZZS9TTvVGNLN8osC4DMf8Pucavo5Sz8yfQJf7qu5C+/9wmM7/g54zJA/LfzthY1YbR90AY5s
awt9Q2tG0x9Ne79h/ivLUcfJa7pvTdLodmwVYn9++WT+KEa8LSDnCw/zOrL8YJoadyPbBGKXoCSu
off36gl5TCzFQ1RSRo21KNYKbBM8EvaWLAL+Kgnb2tkCw/661LF3m73MW88V0c03T9TFn06+E2jS
iHAZMYKAMXCxCDfJGGy2R38h6OOGX25P3nesd8KJz30tUG3NgtQQiEc3m2SoVmdXhKJxl8lDuRkW
qy0sx6f5s54oakxJsHJAsE3rE8Hn+HkXuXMr2VZny+JM7PPoI7Z/jMflKMS3y5eOdaoHrK1X/V7A
+MQ2xVEJIKqELZf9LXYWxbAhfuEAgcsahoOO2GcHviRFcGZIfLI9NO1vwlF2R6wyJNimBZcswZpj
WhQSrF1oasV1T5rOwSf7DFvHWKo6TBeyHju4AjDDKPkTS8It7DTMq4/qgyj9MD9xlR5or3vx1Kp4
juEZIRDO/QvLJ8ppFaQOwbDlg7G1bkc1ZNg72QCi735uTRuuRhED87iia3Kat6Q069qIWDD8hAH4
ftdyQ7zG+uOO9U3v9uJLEjLwW3zg7FcXK4UAnJ7/pM7JEN7n5DyGBs3XPuUckoimvU+th7OnYohJ
yMaT1YYT/adgvwTkIdEiNQ6nvNH4X00wqlhQH5yKNBbazF6W66Pe8OT3q9MR/LhaJ4qlbSXkUOjI
iBrNBjFWg247zijRyxalBF5aE+bi4u+bkVBYicYtNQZiSx/+l7BOjCo5ReE8wJK7GBP/DE6M9pY+
S9yxnKVL+XD5hmWnMFNe9qoDu/dx3tIz62KCxBxcP7sA9Vrg7Q6JY0X7mPyeCrq5ksi/nPsVSBIN
95U8AkBfYosp2UkMvB4msT9RK+n0z6+wG7jaVogzdsnJgnYtgLQjsFvXPAu5nk65i/B6BTdUZzA7
JqIQWQyOSmPlHUvha73qKt9DJXEecCUZ24w8+ogiWrNfBcFczxrfvQagDlVa43npGZdH/gcSBn5I
LwYsuSeuWKIl7hdnu4J+aptTyxf2uKEV1fQU1oOzWeCDQv0ZhSKB9LMvuJy7k/17HDeIakH6BciD
Z1LgNfr5JJW+SXCzU6WYtdP8wP3f0IpFvpH9PpWBPa2/aOeUNUIgEhMrwHWbh8bya0T1n4fGBwR2
9UGgRaMKIYkQ1xxl33cYqqdDhDQSFegdnnK0Fgvs7X7SOhasNDafzkeKkMRR8iOUK+C7S9cIHwLr
E9RAfhjbffLDb1+GCJSKuVCNC3We3jLGq6beYkfujtAjfXjbRX/uC/E55Rbc1Z9SBDWD2JRspY3/
lLJDf8n7xAaamA+O5PAwmM6SgoFh90l/Iz3bTZFxiTDUNE7ZGQKZFgZgR0HmJpHKREBNxBUfqLdL
rpIwfkq/qaRZH/bsB3iYk+HuM0O1Hdr0dEM2F4yPBC3ngFRLUgo2ByjExSQ1anqHmXBEUQr6YsVj
DVFhUbGHB5zM6POxknly4fcqfKD3ZJEs5Ml/ZEGPDOWJxVEbtbTZk+wanZnw+aO+3aT6almRWZ9K
iuhd9rcygDaBgKoZXwDwmMEhZQdAB7SdatvyrYuaC8KADp6J8oBNuKP4R4KLFt8toLHLHmm2OoJl
p2strD2zfJZ9wyphpdcJRLU0MiGVJtCXjBxlMqk4HYxiSqAFB49Q2Zw9O37e8hTYvXfN2NFpDx+g
asoOwh+aETwDXlqH2HKOD16nKzS6ZoFxl2qeKyaVdQ1ujA/HTppiFHMEBFyXdRjc9I+yhBc/i6QC
EoHz7I4oIUdhnrhgIyrt5ELeMj897mLKG2lqiIH1qaiOnwPH4JU1LpzItgUVbTPYCNbEWVID+1G8
WzXdFiVHF9v+Z6w/amJVhtJfxtifPGVJHjyOWBfjM42znr1N8KfuKXzWRnPHOwpJOQgNx09MxxEP
DeXD8Bsay52FXxCypdMtPo4WVK6+Eta40mtOIveG95FzRdnxAaLoJJK2Sy7yB8g6KtTfXzV+GO26
xwe8nUAeP3Vz1T5SCRSN69XIzWfmbOAmtrBaC7PGdPCSOTKZUAqpzh72szSYvEM0OVPCHKiO/hwl
MLrlkhILA+mX2rS/DqQI62vOLq3qgJhmSYVGe1kHqzITgACq5EVfQX1qzwBYwqlTcOYGV9Gta4nn
tGVLtsW/RCUyD2uJifRF5bLNjtV1gtdaVm+xnS7Ai8SEo09n5PoipzLSQbUARMRV6fyX4mP2ZkdY
e9nJ5tkqcu8OP0TcKVOsrH+rCoONVsWHshN5d5PVMkTyCp+xZeDKRFkXkeGVL3G+nd6ESyUCYoGu
62gcIhWP7JMPfMiYB0JgVW6km10Kh1tu+2gFzWVQCxQm3rIaK1IoaJezIhIk2TA9FSGolDMJXZ49
APl461cywmkQ+cEdwo63pwgpLWFPXBvzk22Xl6zeg3EOU/uk3VwvRJbM4EhzxKXAYSadGd2WKt7i
M8YCJYWiL5rdKBfRB+KsLVoJeJRhEh1cmYQPQqHnifUuGDXJT9U9DX5zDvVelDdZH3HpXZhxAm4d
X0jXN7n3w5H3knyo7Emlq2LFX69x9wjosl/EHDy/BoVJ3vJaSrGhlZMkK1PxDbSJLneGjkKr7YFo
cZefo3aTeNgHA3RE1p39SlQTDGQgsqt54jJrCjqredahBBstrlKohUKukZ0EwAqvfMVxzwso1We7
I3qiJkfyCZUOfYGM57CSEFHpCPeoesnytzEId6H/EtRFkuMZosO/cywRgHXIKpl8FJR4NENGLBYL
SzeHprKHbD/XyxW5FROQnqcSak72fERsP2xx9ye3KNK4n2fAro2A71F35mhoAvxXcXsE04/a0Mvs
cGIDi7DiLHWro2bVDr3czOir/ftQAQDt6g9Jgh8I2dCWXKJWm9QdSI8Vvz13uwtfkzfC1kwD/Dsu
VWqHMcJ/+z1t7op5UnuoqTRX6LhvpQkgMBQNb431d0fDQypxWqNlRyYuuB4a8aqD/BGMQN9wis6k
XXyosqTFdnEVjU2BTglNsF2KmH23aFvJL+h1XbOjcB37NIWA4tGtQGseGXeNnqvYcutH/8783col
RzU2oqwRXO99rTraXQzlJJrZ5Di6zWh0yFzvtNN/bi8VVVHJQo6Nv89pdjdLmwWJ5jDk34O0SPPQ
zxAk6f/Qmki+e4nPHSfq5mbx0gHUfnqv58IH5T47tgG4L0/RCmb3wATROi7d1ceOX8mmkjyVo1LF
9Kb1L+SUPCLC9JTvOJYhefIh88wqRA0QyThDC5oOPXI6iRiLHNp2cJV6fX8o80K+Vxbds1owqPuF
yi9bo1DCk80RegF2Q/JVDFigt0oeSAHVYvfXVnHvlXujx+lBlyCGmpN3dkZBe6LD4Y072erpSHAZ
x9YuDi2ado2Lsrl7L/DN2uqE7SzeOWLQDrbBBXs8FkXJdYUp5fpS72+ztP/NctWbvKEb/qYXRXh8
iIcN5l92YzYY5zlAwN5/a152NQQXF2OhTGvX6x8vrfuYN0PyXoBiPdQyhtxULypXVb30WD5Ce9MC
XXigLxHgZesJ7WFMqv3Ww+bX3ueYoZ+Gtv229e625sNKcxKLiZRjQhTW0iScV03+FX6PEx6GaWKS
aXthlbtm+Il8HD2FL7tZYzVbFyNIJgncBquLseD9oNiz1sogm1OCydGgDgmXgJeYzlJFv3nHGcZf
EscfIq+UBwmhP3byPyg7EWmJUoXohpUdvIXSasnl5uXOXSspsi5iSTaPIFXRm4XoW24Vr5HTBK+y
UERP5savUy6Cr/P5YjBGxhESfKEbAAIjCJrZQfyTfRlNwgNo7dsHKH1XNUB1QqDgk7pAC7xjE6pt
C/f7GQ45lbJx6KO3EKdjkDGQrmYVdkbJwMyftpqQg5ywiIzPq29mi9g+baPa1y9roOXfYUFKzVa7
GJtiUGC3LQz9jRrDD5q0A4ajKnFk8N7/rwqN3UeVmUJxo7s9EboEVnzpjVep4TAruPKo4VXWt4ud
N5p5dLE7xzM4oouVW/q+wWLrzQw1u4Rj2jX7Mkf9gbjOvAM9gFOlr04nodeeL4pocVXa4+S+07/W
rXv0o54nnZoXrG5EROyl03n+vqvU8Xc/PJIoTy609MsczhzTBC2KshKQIyRu5RlnmEsW4FXBRUZe
ah7zgOZYLyMR9IZLueuJPN4kQ16wuUY6/EL7EY7h+aRKnQVdi15ZS7SLPx8gQ7VQh1U5SZWul7lb
nmAUJpfohkcKiwb75FJXuIJvHZ8I097DP9sh594g+mbZ9OBpJwSHoaxQorDhGhEL5LL4F3L3V0Lv
xiSwvB2tPH75QfWzzRbkQ56+wRVYQItHbaKYsjm8KIKwnHfqX3L0gqhu90fmgQ4ylhqBWJQUeIUc
I2sj5LxgFE7AMoo7BPR9Nmcz/wyevy23a9BPs4g+82gYbu8FTLC6OQ89NWXGUbh4K/F6pdLKZjKF
kpueAIduI/m/gmxb0TwTSII3q4G/+3Y5EPVCxNGz1+2oPdLsYnmIuZessaVOTjqdAtxJ1G8qtNCZ
crsC1AxJwvZUpCvwfcWJHx5rTw9mm88jTwlugEDE8Jio8U5TcYBHBAl8RRTc63gVh8NPuig/npOx
I+4fE1NCawoP1INtfqw2VJrn5KBx9U4sDzqZnKUyuUV3uQotOWJjgawYaGmlB/6zpzu03xIlL25U
HEqxIaDlX7gYM191jLiUJ6GHpgt7cRzxvXdFo3eYv0qnj5rxLSurrBivDtaFXTnXfQ1OnFBHa6Vl
kwah/+KSyve3LUOO8uyeQNQTBsnIMWo3XTlh/3o8Dw+gi+xVlECiUrHMr9mRo4HJSHrd3MgGOsw7
mMf4JeHRLa/pmTYBL70pmdEBbL2WUtj296k12nijoXFWrlgck4GXYz4/0yZ5kIiGXqfuB+yrXmf/
xCeNVWqtTiQWviAD8mh8vFInecolUVxJ0yZjEaqVdtNnbmr3Kh2GsxmcqKlOgSp0Io44eWsAb3ie
XphJe3X83po3uXZjg0ywZuKgpK8cf31+HzQDdRAU0jXDMVEPtzK8cZOrFDGShq/B2gIuct95PtTc
2ftfRmYmu/oEDUQAE8MvTyLmDRmdyH88sfgvJQlceAFupZtfoZpuoti7SbAKyTv2oaIXcYtWCXdh
0kYaM2W3ropE688rFokqSp6nqWhk02ylLPRpDKSD23ZJp3j+DAYnN0CwtP9gheaAk85nQ0A3FSSi
cYHlnYq8JXEIpUERiSaoywdjvO96gYm6FnErHVY3VPXnsPqMncPr7ifbskaTdPGsoFDGIa2gpWp0
5nme4MOGS4LrzZarISbNCkbLpa/kOjG7sx+jPGzH0+xLMPCyQI+GU4rbFiW+seWTAjrREWCQbVh3
fFro+SvS3ekd1NdoB4+o1QpYBuuZw5xzNAsCm7SAls/T0LsPYP2bzF4GDHCzcLfB//gbZAAhvkmk
q+WUSWUwnIxwJS97onQasg71OPadnMPuQWCcKNkpZyLfMPC6hb6OjuonJjmQekBQWuDMJ3Kp1hUu
6McaHr+DVYaw4tSWXIKK1mSkAYYjqxmWTOgrJBgENeGP8Iavdxehvhmlw7xEy2lcpcZ67l2eAt7D
wN0aH2lGGG27Oa17MBstS3dUcgkIR+eP2xjW9kE/QrQZWBz03yVMQ+ZQXtFaMkivAv+LkUufu+6w
qUOziPWkB1bWmStt1f8zPAJKKJ6mcA6s1vCeLoxKY4DOCcFBHLk8dQwaK6OV446O0mApBreJqc1D
wwwRLNTmWeovFtE+izPK6edfGPI/MZkFR6uueK+GXTkjkvi53pAFqR5qLmjJytDwhFSCQ3smIUNS
LMNA3+/KcqfxvqtHgDT4wfp0rEfsYfkcpvXiFA84ujx9B1rLTlYxgQLOiaXnjNWmfR/wC/F2swPi
+rfyCkHLNtED6F5u8GIkE8+D5M1xB7t6/SFuxnk0FEXz3IcyRFjKwrAkQRyBoAHCYZGwG9t9s2w5
xwrh06lThnd5XGbUDTfXuIE/ZgUBPjOMomGFRpnEEQ7Q6yiWtPwYB4zRdPV1q/WC9yzbPaQKfbQG
vyZfP2ci67dDbQFgllp1M57S3QFAzhYyniLbzgYexP1thnl4z17WM0XrX0Ar9nrLX6UQqYysH8xK
xJ+ibl2VIcSfuqTupu8GEBi4p2FPAPbJspr9V2+ofnVmRK1tZAvAq09g0N0pJkGIN8tKjZxhtItl
HBJhG9EvGNPwN1n9gBPEsm0JXV9Y79BfPVZ266Z2K7fkkzUg8sB8XnVstQ4G980NVcRJNCwAFoQ/
4yNoNQUwfzTd+DxxkJPUWucY7nsXtH+tOxO96Z8VJwFAoNJk1ZorwcxV5HLuxUAQo1RvVZwHkxzw
utnaM8pwDU+SgvKQA1CmWucnzjJm2v8HIRK0L4L4uzp+Yv/JXfVHcvxeR3xJIQcXCXr5033v5ybj
UfxcYJ287XFTrRCMjyeN4V7PJ3ocGK9sLNmOTupzanhnKa+fSEizWm5Lxu6eW9t1hEGZ4vAzR3Q3
RPG4Ligne0eRSEzAbm1pthLw60oBqDee5IeN7J3b39SeDyutfOfzv+Dk3SFdhoHt3/GZKoQanxmw
+YTQ8Wt/pEflxf3ew+mJ6i/hCbzwd+tLS2ZxncZsFGqF3x87mJFqI0Sva4ZBftuUYZLEoRqRkCLX
PF4QAIO/Ln5eswg1Q1rJfofQWk1RuqqP3+AHnYLfQB+BjlX/0x/PxmPYHxiP3RYOlHuEBwsEFzFK
JAjmzlkYPXsadLhkxmqzPhn3V3cjT7s0ABATLxbNUy8cc9I19ZFPvURj7HkZRIxr3rCIYJ3pe0z2
GhlsZvgXDE6Dic6NfzkJVvVieCu71rAImewVl1vbunX6YV/bORc3/t5aM5m9qARJfk5Yi2ygUGAJ
F0QhCF/uIrLKAPYEC/dtGz5aiffZAZjmZkT7RyMLeTKqdXWvOGPHG338R4r//vPVNQgpbXXi6r5Y
aJ/fnYQ1W38Yu8X69r3w/yERt6ogYapfC8SmVMpGPtkywviBUa/g/CuwDRIfhxfR9EPG4hd0jDGG
EBPehwYcTW91y9MWRu0tODK255zeWdLdHn0Fw7ugCvz0lrL7armEoSLGRxQIuVcfD8KLr8hyF6fs
pddhtH20A95xeJjporYg0TYDsINi4dU/7TEWkJfp8foZA4gIiUGQB73Soa8s/1N0gPegzrppDxYC
zc7fdYnRj8puRymbdfCgC+EYg8N8HlEtriP5HoRN8chdgfwkG+hMSH74BsVxOErFVllonxcwSJyL
YkNKAQGa2fqx+K0A3TI2Q3/YKXngm1XO/m+p8XlCgRfngiakmOPmCErjwuXhu9kV3NYJ+LZqVHOe
MUP0Jq4UmRxVqoOE9Wkt7PZzxXUAN5hsUIjknk4GH9wjAOGOL2+GoBk+3vlqQ30Ae+JT0idw+RiB
LFSUVt7qmQWTtQl2u5BlARxfKmRWzGsqGybksh1TjWvYW6LEsXjMSmw4T4+KCAurpHXlI4eAOR40
54PSH/DF0mwuWdVaQE90XU1bHrI//kTs/9v0QLnTYo/DmxAQS5ErmIETbOiIxb4tam1n9MxGydiF
Q/KnuSdiwrMHz/xUE7qRaDP/ax5bxhZO7VHAFeUK+/C9i+K/IPVoYZBMB+lnZ2lluywp5MIGhHJM
tBJZ1+EB+VNGBmx5phwH8Bx1Hx9fnYXGGqeQ4CDxp9SY5Fg2zkWzqGOJowXgVjbk+S98qqJ1736L
aZz93GbIbt0Lmnd2skM98D1DhMFkxRUVRnR+tJLUQ5LBFjR+SHlMuXCvXVooT+8tty0VvaIXwfrn
5xKSpelOloXwOWOPmNCyrzHvUUCZz9MvFGNW8G6MqV7yl2QXiC7fsg+5N5OsNHcuw1WpdEWQMtv+
TwxPxOGNek7H9/WToaEWESQoDVYtC0uxs82xP8AUii7E2QH4OjVMKxPN6nc7K4kkM255BxylN7y/
jsDeDbiILh+To8k7segjLuMzJOM0O2n5F7nhAxSRcM2GfHhAlLdjSLgYENWR2uDJht8jBMFFhrS0
EM6fey98VzQ4eKKFAnd5Klt/PpojA0YEzAag+pnb+1WtGKLtNS6SHgOTOgjulca7mrxu+/bYjE9v
2iuPDpwfIRaic8SEdX8yGFwWMx/SL1LpgpqQ2wR9znJ2skWBIErFNqT3m75nG0jWJzVHoGl7JaJ3
ONfSbAQifcVGf+XW15ICvNL80Ujw/kbBheizFKdnHjmqQAxEPhSz3rmMtU3C0ktnnOZe6uF1reUN
1200ZbBdosn8WzaFDR1CJF/sboWfkiwxPTtieX20/0/8Q6pB6AhBmZCchXU516KBD6P+tTGm4FD4
Y0LQQv7ZeUWxaeaBBz4rTzzqtxnvQ0mLsTJbvRlCs/JQGIB+D22OjW7iJpUIJOL6NGqecCdE0O2M
WC+9kEvUzag/YlaXKmAyHIpgjtKWb5DnKIPJw6a0j6jKIIyCsPrf7ar0kD8PCJ/DF0Yk1glFlBXQ
VD+P6xox1/Wez875Al7dWRsF5jrKmGZoTga+SD8gX7CI9nYEJsZ+sifZ1kqk6R8E0nkkkWmj+2U3
qNSso2qYgymt4YCWSAb3bGpDUu1EfN/SQ78FD4b1RY9cb7oXczvlPE9EVdngEN6LL/yInvLdGQb+
f9upAQ7Wu/mzm8OrkPkQdVR9lJkyYF9Z78+cYoh+RbVfTQNKe7mc+7M5KOnq0+Y888SAZ61hjVyt
RJ1Btrwe+z4Iq26onQs8thjsaDEqeqxIwxa+40JGp1HiOGFoQmCxVwhls5YFQ6cfBYwPJvry2+L5
dwUViMm3Fp03xNxrqdMqrc21awomKBfQrgXSYJmiCGWnLmVBGw7xBRq7qv7PM4ZilKR1rLXNqNR5
TNoYEwcU79fl4d5a0rSet9hR8uqYgtgeuno3jURybtUEo7PRCPq/pmNKjW6a9O2V35t7Wn7eTMjb
jinSn5hUe51BKt3dZeqve8oT0QOrL7NCEz3ApwU36SlmLPMdEDM6Ab+ap3lPU9obl6KxYASPu1Ya
bKouaqjEB3Kr45RhOsqx0gaXANTCh8GvznhrJIGtjmzo/5QaV6CKWUORxAv+FS323H1RlZOJNBa5
crXgnnRXfGSmtulbOftJVpPKhQLZo9rB3UZofQXNiNN2+qwiUbopr24cJ8322ebNZlaY7fCOnqQn
211yIjB2WcrU8jrLAsyNmwuFM1ytEHPvpodIFLVggmEQ5EHPBDr68eoMrfV0qiI6G/556AyLNhgQ
6yI6LuUdbjWPxGG80mB9YVfKmJNRX1ow9cYzTufKH9d9Ux2n6OAyB7KxjX+rlQJNTmgIGCengvee
wmrrbaY41nvHMvP43WBX1u5Dsbr51Z//Tzwa+dhRPw+JLEUKLl9ClpmAqgMcAR2SUUmwQupcG4th
3bkGV1IcSYvMbXCaygKKoHisXjMlfcLcU0bOUJH8Wl/17+iXQ+rzdyIjVWuHWrb6X8bcjXT608eW
ejsISAGJL9KXZ+4wDYpmepP7yBcnNslGWmaGeexzB1n5ExRsJgfM+6vwdQNq13fj41CHzeuuGXbu
oksuRkODQPUjj75cmrtxt1d6fL0vQOKRVbWihTpnQUwKNFbcrYGb5CzSViIuHu0fQTWa0VquqtD4
ioTUX19llyANlsFe7ylTK6sI70Y2rLSnYvJ6NQX3MgIzQ6BR3sjpAYmEWUPvY4N3VrbjcC0VkCNO
2XMbG8pjNBGoVuOwW+/IUDl2wIPfMy0lxPX2JTO2CNX8kBRPuVFhf/AdFgZD8gNN89hIJeDA6V2D
47emb3Xfaurcj1/IJU2OVJncBGdDvLFeP4FxfZ7AXaJR0QYsE4p3l9TRkQUAB/hWFAhuF6BNPx/7
kpgyH0LZJLKF/C8YNWhKBcbChntXOzFIsym99rCQkoXzM/AuoCOUHY+3hn0dNJ00hJDICesvXfTC
9f5G/aY56/KssBRaC/EsBZTzO0cygUhw8dDk/5DKgM+/fwiR5kbhfctsJpqxc/5BvxYKRLnZOzwK
woblEc0QewFG831txazJouhMgzW2Z4f/fsvmb/sITWh80zxAGrM5uP6Ux3/qKg0oh21ZhIDwUO1o
25U31Njl/XSf7C1hOc8TiQd3wZFBIbhUvwJ+LxYgbF5DuchWk4iwfpchEuEkjgiUMPH7TmeDWhvr
zN9AxM0bua9hLXjF
`protect end_protected
