-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GZfFTU+fZDVm/lbtzKmrvsGBiJB3sysKs1ue27FLJbc/SyWwjy9pBOZCly/3+kB0J2V34FPkQxL6
vp3l0Qw2ISNOcg3gmB9lPHEPiNWS6Li+IqnrRRXhSvaTuyEHwlBFRkWok84+JUrH/VUcYeMYn4ui
fwm3fjfn98kh/4h+xo020MIZqAAt/liPVPjoseYNNVqZ90PCBWwDBmcbBfKLqlKnKP2+02T1DphJ
ev0MithGJXjd+BPTnpSb5dkMGXFmRj+rNP4vIFeF4G7EXYaCxgtbcb7SDA0/Nec3PDmDcV6TPAPw
5dONnbz1pT1B2vcnDWOTYZLtwUoeEOkiDDLIqQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5168)
`protect data_block
Sl8VDu86uCN+LqPqlyUJswrMhdPozKEhCCCk0SbLjD//hvAKNtly856qRXIhBQTM/fVU+IZE6hlx
6OQxN3iuOx25URFHeecynlV2tbxgx6fAZDnkUQizyERwAdxmGbA0atn7YL6pX5x3cr0j8e6Px0lr
ydAiLdhYBeczvqYb76FLVE2YIBMxoIW+XDflY3hHiUGGCqC/BGd5kNxJI1C9MSgOrnWxXxiVnuU+
MKflQxN4LRJ3Hp+c/+2QzyRdEWIO9OEg3uxckqCZKnTTapWA/ykLWT+c52d2HmK/DBHsUUZMEeyl
azHNO61x6Nd4eOHPm8ND3L6IMkId2yy3mNpDs7Zt/CvP2uO0ERQLDt3iSVkqqP2ySpvM0pxf/245
2FuIPz8AbpjFkHnl6ne3hjHpf0Q0wZS6kOBjN9dgD9t+cY9JBSxMy77r19hdA86e5Y5deFBdDalu
bgbf/12N+ZVNqb3s6oFQZQmWDrPiy4l4aD47NDbxhrNr6HfKpjCed5EPTqOiSZhFrl0R4UMjtRoX
yXLVEjH/fv5pZyXcCY/coMuN2BsRsTmWqDMLHDCM5aoY7Q8cLgQnSke3YfVOdvHR8l22+IL6Naco
BRUlbgXVDMpfJ4ZfTwFM2VzemGM6PgXQAaNiacTh+GLFCX8EYY9O1xC3xGsXaZCS3LYBRmXa8OOK
r4ONGOoSt7jTAf15SKHqDtaMH/2+yyCHAkerm4BF+9lpKqKIs3QQJXqsylMFTh8ra4CZSyl5lpFi
485tbgszaCO+xYy3l3yTaIOOFqFqWVl46u4JNfSs5iwufduVZUMSYtm7Fdc63mW6XJZ/Bvp9w5Cv
kithK5TsDUR50C+QwA7XywvMf5aHNL7Aa0PLNZlWwPRSPU1zoOfN5X+DvD2DsyNq2uqZFeFGcnzD
7YQo2P+zoh6fBLphhrmIpriqD+fGJXVQnlEv/m6UESirzo5b3BcnbnocXhivi+65DJdl2Yg3ansL
5lsg21UayCk3hD3TGbROBy8lXwTsLt7/TVd3K9WQcEozgxvsWkuamb73mnD6RZRkPD7EgFLk2gKG
k9XXgA+81FNWz1JMgL9xn/Q1Ncj7axg6e2DI6hjvp+UdVpSsnE/jv14FMn4tfJUyQ8HVVjQOetbk
KGEzEG7/zlSBqJv2mqEDCgqlYiAtM0OWcNMCU9v0zvP1uw/9tCqQW6PAlMN12NrIs+JeOxUNU/WV
bmHPW5uRmn6/acANvU9GtJCTmGdpG5A5WBw33Av9384iI3Uq+JIGdlmJ1lnzDvf3sKUPt9xzWMgl
JaCXr43yTrH7oJLVaqXmXWwfpQInKvFXWrQL1xccQKgdza94pgr8aZxcQEsq7W3r7GhENV74ZQ64
EF/UmU1roBQ0kTSsfaxc3HpheRspVCSKENtXXpoFQGjH6NHYOS4orMw+yhzuLA5CnRqinieiVfNR
V+TG9W82cs//VqzF0Mxt7A6z2l9zZhNYYJbTla29tS9afaTYrb9oW4fDGYIAORHPJNAPnqBY1btZ
P4taClBo4400mz8dePcQzNniZc5zOMbJ4VDMMR3c3Q9uKMPc5XH8W6S67FyopDRwgji44koIAiv8
PKKicGR4Re3e5vInY3Krdn/V267tCx6ExffLk4TZdzVAIyHEXdjBvE2tv8CNwwkThHKpSrvraXdU
Wk3ghTMQ1LjTOE8F7KM71N0Vo6gn2EkcwSSC4tE1xt/roKooBbQrpMRc/6T2s+efhXs/GnazOm9F
WZadUin0eSg1vYrCS0rdawJa1BV7si5b2feVUbB9kAMMRJo420AupgPS0cCTFRYGJK0/GlwG0YvO
se3XROzPPNQRR9i2nAKgFV965eAcgHdPde1GsmtgSAx1KvHvDBL7/0HPoyO76LCtJ0sGLSXypZtZ
42e2QSID9obLrtx7cZZwSWGjA+7PEnE7+5LU7MYU1hFWbIEbYu+mkGYDRistqUTEyfTAYFRQMKFX
gauqgjKXTRhujdN/Ek3MxAymr+ZsxqkhHOv85tazGIydkXD7661SH7bnodMn0mQKVCXzQQLVOWtU
V/h1eYre5Y5n2+PIShOwnJMJJTy+ZiET4CKMnuxVmVIux/170qsDFQLMisUF/G0SYEeJSzifobzQ
CURaWhTmjOTqRc96ug8XvZF7oyNXd8OWhWCRcJo0G0sZQVWwtcfXXhwt9LnMowg8sHsDD5stitYb
1DCsp4HnnQT62v8tPlaiipWnrjzEUSGcd6lhmE7LFZtmZp3N9K9OkVUSUvtTEh9m5UO3uH6njhpP
gVaOnpiFEsKGgcObpwyKkZ6joafgRP4BUafL7dCj1OBiQh5igvI4SScuJ0Oemr/RD83MTXgMlnrg
XW68ez0JCH6AfbUlIzY2BS1/t2JzwPoHcINjxYrx0FZGBoH5UPb9kgn4czl70py7IW9KxRag+yqe
UoBEu+VgQvLgl/5j7vU2IzM+cZQoUQVDQovtZKif9szzHryhllUAqQhGxQ58DRvckAhMtFVwO2it
29lL0sBrZEj9s/JCy14ljuv7MlUFuQ6otN70jXd+yD+n/w4GSdAmGANVnggdXhEP58UDYS2bHFxC
qTYT4IBr6VFzDpq5x1IOvMxDBJduPHMGOJ32TFV8WxMShm8VkzlZ+C1w2GAt2NZWlmjsdtvkIL1I
9WZTMGCOpSMQbLQSzfwMWs+6MeJprMEoMBhIJldIUccZqjdk5aXiIFeznkOtAUWdzrLQaX7sENBF
aAzVEP3+qMU5gMHZh4fLcSEvBn4B7beTWCzPN9A0WO+D9G2kZIS/NHLTDXdHK5Ftt4mUNV5DpFxH
cz5dSlge+fBiUNPsx5zUyOR6U0u/X9H3pi2OMxixBV+9ua6uiGPuRKEPXipaZmclWSkbruu7F9f1
vKJYI9P0LcJBGvxnvE+rM9mOvDzJnZGhyYWKqg5aS0TEOpXKYZzhwjGBzXEInYkW6q3ivSdo6WRT
kZ3YLlzed0nPArguVXI9flUj5JcPf1C8SqBpMSTTbxRx+6mZjU3LcqudFVsHOssg2kJbN2x2vdCn
aCrGnsW1ZFpF1Ey9Uzrr0ox4rK9y5zo3YnzodA4nWi0N10mJPCYjo8tOACc2lvKiT9D1S2zd/Nk0
I5ZLlIjmQLrLZZiLwDp2FjaQ77JpbP3U7tfJSWL+c73PZvKILltfUqDBL2ewrKhjxZRULmFWoAcm
Kt96MekAxBPtRRPnV3VyTzbRmwzwV1KNLJ4JAgzylVAp7bAGLxkZ0n1hgaIpvrOUw4BGi14vNuXC
+TIUxR8CXTBmQ/xfcJWgd8TjX9vXTVGNtmEXXLqaIqZTBJN9VDIRc7B3PUNNZOpzpLjcmtKm5tnP
B5nsSplkPV5dNtajzc9zV/a0zNckhA5vqv/dNF1Lf4hJhnvlOger0JQU3wMic3MfVCYUl+6/U1vC
f3RwAzgAJUUzJ4OJDs392IUcmCF1jH06www/+M6cGb31XtY02evaf9/nuDHPAMTVZPYtW6cjTXpb
bpZ1jpOleyvArbwoyrjqBXg8miMOLOpBjIFY3loICcb0yr46h7vZLBXHRaZkq53TjJxv3h0VgYsI
ux4QPRaMWAuXz8bTrmnl2rnaE9aJ1NuUvQTv6vvWwChYYVYm1HD8pHoxxDi4Y52P9PEiS6fARQPc
pgn9ckopXjeYQ6PosTFG3+pX86TTGcNthKIXXuV2kxo3yDt64T/vZAjwwbYtqMOVQ8gMG0y1nEMO
HsomgWQ6uCdQNY9iHFNKeOMNO7oSwOjRUo7Qecg8dXCIhdO2lTs4t4kA250H06ANua5XDI+pkNfg
NcdxC0Ztm1Uw37JN8IjUlLGJu+EwuGU1FeqPj8UQN7ELGhyuBjSwmSEZi6aEzGuAUNk6YeuZD1ww
nU+U9pAx0REXiCPz/RVloAYb5jVfh35c7cVd3bQ3O8OaV0n/NjL6CreFLRIxHzsfbubsiMerBe9N
ocCeuqONvI+8DJiJRQoUxaFmXG+BjJzy/IP5MfGmt7JZ1QUuj5NDmGra0uqbg8l43dRME5V2/LF4
gdW9tWXYWEQ9r1uC/KHl0YKOSSDVaj66uVTSinQuFOgydcXhteOd2DXS8OjHTWMcZIbnNSAMRtaw
SiGfKFs8rIiXP2S1dhOAdU2daRkEfErotN9H5WBIUu2A78zWFfZpMGA5iRosZSuMc90M5VjPqfZn
L8dS3qa+J8XGOYPQUb0ZAVOPiQxUMFkbSOnG0qaEf1ayklFd0EThEgr3VgEwix49mVuXt0e+TIzj
EICQTWB3q+1nf1QMaX0JbXlSzpy76uUVl5t0H4+34OR16w2WCRm0Sf7SJiGXN5iEdah0rKlF7KdQ
5DHfDPZldMzligXYLMofvaQA5I2J1JnxcQhmNAV52LWUi+K0mM3/inluUYlIPM+BHsr20nK+MuLS
NjBORwfpN1qpT3xKvdj28XfVNtOh/xAdlzJNnzWkHgXcPubffhJuo8cnDxq6lWGx88INvXk4yNlV
dpLRDFZrcnk2nUJtsR8d4rsdB1q32KruZ/37UdRPftliuvSHihHMOCRIJGhQtO4DUWmY/8CNaUzr
DmI7j8A2AZkkRndyrAWS8XRMi9M945vDaL9nsBMOg1buY8xNomrrIozw0yAK5hEZEkV6o+9YPANB
0rv/cPB+mUwX4FZvEuGSVx+mAqvt6Xek1X7Jm1ubQ5dfTA74bWyKOG+bTgMT28jD59AR/kCFUN5s
7dunY/rtWXe/O8yXVg8O85sxYTR3lYA7w4/bb56f+Czf+AUxPRejs7NsDOuXpYu1csJjq+wz61yi
/lmwQ9k9NGjKfHlvNY4O7TBFjNyvLnGbHT+nmCIMaoXU6xl97VBQW3YQtu8SEvncjj2gW9WENZlc
5VPM9n0aPwbO/tDr0W3SudZ9seDvBTxbjJoI9j0BYe2ftf16EVxdGD3jmnTbi1rS4+haOKvhTeL4
DHTdha81KNiqBFGzgf085eIRFkRfM3uI7BQO0g4ZU+WmNlEqaM3w+uXd9utqa8Tx5jSgJDt4SIDI
4IYQpcaD8g1+wYiImsffrTtZ4if6Xf78iCkZcrKvqtjC8H8gYreUvSd4vnlY9wWqHOVFpwpfz9vh
i4ceXkx2/1QFqpsVdx13eciE41FlawZUqqkBW195PwE1Mx6ed/v2u+PWauCoFAX24wKS1DOp8KEI
SIfpYoQaQQgNoneauOT1LXroxr4/pAJWxkBk3edpBVeet9p8j8IoHHvk6Tk01ZBvxuKVx8khg/Gg
h8sgbNc0qb40aMNfbqKMlJVp181aPIZPoL17BA9rxvgFm9Mt/awGL9FH45rJMQeijX9HdfZOoHIT
OV5pYkvChTkwl4ebqQl9/4SIH23/HxcP1YJVH2Vl9dYouLaBXqx+KCIQULaHkAdaJU18gO0CRv5G
7bqjUp6kVC/yaQu+FwDQjFkLziORgvqfGFhZz2SAIbMojeg7tvofvKNIOhpyFenn6RpWjkUaBsli
S6ENxcHwwOR72ONV7lSHYflGowg+GUX+ofSj6d52k+C1kVSBfInUroaK27Q9a4BrfqVPrtdX68ni
2YaIqJswnkjBen68FNloUQyZWVuhrbvQM6XnbrR1PVX+hgXIk8Pfa2K9U/mgMVD16hbldlfDBhRv
NWZ14dmeHpY9WTJArFJ3WSrXFUH4GoFIPYTT2qLQB+RtghojRnn1T+k91/f5vSp11UAdUsz27guL
RCvZ5fw5Cb2Bx0ojKWA5BI2YfPfEOLcJzbqF8/7Y7sT/IxDftMp5dPdV5lMPdFmz1wF5irR3nHPN
IAQw6akgsOQD+2l53/HHyauacILiQ8a7KmPOUK4Yer2n0CdjVflmXgieYiUiJRb+DYwcz7/b3hGM
bcdXjdgs3OAvJ5IGp2ZGUNKlUODKYTAD+XgDjeIL+Ds+Vyn37XygHPk5VR40srX/Pni42OKR8gHu
hGHRq3nU0wcSReXGdXHt36iyO0TjaAd2QJd/5CGQqMTEO1Le0XaP+DkF00RcCPy6cjrzL8m/DMZf
XyVNeZmlWJQDaoAYcrIG3tTUQpoSDJ0gSF3HxqA/0VOH9qx75gqAIynrFvnHBxdvTgrCHe+lOsiu
UwnB4OlFakjiERcW+pJvU2aWv5109Qy6r8QBEdawzdCxnDuBF61brgi9X2ve1YP21J4vMq9KZCtS
lpR3EHXsT9CVmtWuGmF60jmjV6LbAAqIz3uoBk4/TqSxJvo7CEfI4Zao7R601ZsNaBGGJDFcKfYL
XcwSDzy1ye83M4sc/3OZMVo3vuinqgmTQBki9XUvYrBPqGmTYlL4lU7h18GbnKXfQ4e8SPQsiqj4
MdMYQx1Ub0iLAh/EoXh9B86HYM2dOJ8QWfQOFoYp1nnkRPUuk0oqsrw3ccqHlaacxMbmTe8pJ6v+
1Waybh19CnM1eUPVG1kxKxrTj/z+winapfXSODhevmTfEpYLNj6UjkLx3nS+6uoN2j+UpmJ6XVXX
Mt84xyEJu0ovo/RTIVrr89KVF7/U+3Toi86jZ8GvPwn53q+b/XvPyy9QQZiOjM4eJjzWpOkxUGOR
yMAG6OQkXs/2CixoCP1l62bLp+eHvkU2TWLMQ+V9UbuyupTKrIQldAiAESBhTtiJ+VrPECjCy/Xd
g2yKqyU0p6aMAWQsM3G0Mxa7FzMZpnv4yG4F81GuVmMB+DRMbYm2sn+pMp+Z93+7zs2bRP5wgg6E
HTF5nRYnYhe3Z8DR58i6GqGE3Srb2wXNIjC6yBhij1TRX6uF65U/G1XULxIhNvAoh8YmoZ4Z8sj4
xA29le43MgsurctrWf3RiJGHuQk/Qd+FDQfWTKXDwA4LWQdZZa1rCRgkM1g98/HZTM+0/rQt8Yv4
n5M9PLXbkTVTzHYXGugCyyz6+DNWQ17KxoCpI/At2mtrAUYt0bY=
`protect end_protected
