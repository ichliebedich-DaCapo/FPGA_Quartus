-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZvdIjiI/GZzD8+hO58ls6iSTwG73tkXhrU5X47b1EdS8VBWVLP2eoWSohYt/lXfeGFg3SWf7SP0k
NxZurDjWOuEBETwI2wnyCITevuV+FVCQu7UXvBhHtm8QIuWaYTB0gGAv0HsS68tX4eKnYLZO8t5N
CKi1Hk+si6cJ8wNm+HMwxRac+ZAowGJ1FINyUXIc6IUFTjwNMKqeceL/T5nbcIJ+neeK+4Mo1wgP
FtX0fRJ+pZSTysC9cxaXiRZuMbB+2HWpMx2r0O0P+qFBGSNLGI68P7GYEiGSLFGs2mLG9E+NlNgq
HZBH9bt7SPZ5HU9AkMYlAZxzW9r0HN5LGRDrLg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37232)
`protect data_block
NwnbqsLiz0fpXnsAWR4nBy+rcwxOUs75EASIMoB/80j2mQLjtpmNelRT7g6s9bmyWqpJiF9JLKXr
xpsNLljXCtROA8grwdo72tlJ/swpp73s3W9S8fnKMKHbGnDtoPOvfhWc+DV7zCI6nhNYFrtPQdYt
583gmImxkY/w5lDOcrdvHVk0tEOpWPPfeN5Ha0Zvxe0GiRvJFlWrzgU+7h0WHlmIcZC8X4U6Vb+o
X7VMeIof958EfN7ATFRzWncSAtoUL3L6H3pfA9FSmcJXPxgjTHZ+y4MeKzFDEEtZc6tFn+gGrvTM
BEysnTUhlOFRac5NzwnLG4hlERf//OEvmOP2DtYo/BiaFTmKWcPkSFNdN1xrmwM/JNS7tUjnXMnd
sg8TNoqbzJG4rO8lDXUATjv9qVUGRqU61oQfWf/y/42PI845I+h4FrwJJO1ndKa3dLyk8pUTHFI3
ev6aBq3xrLpMnkuS8svIBmztKGpEmqE4bW93fhACn5KTqsFXVUsTwGpLo+jIMSkA49JS8J1btGEz
tmnUlJhvQ7iA9+Melyiwey+pUXYMvjd9e/8eAfNqnWSfM+gWwRpekBESe7Ya9VX9yu/bKf2Ta2Hd
KU4dUlEE2X4lUZ9oBu+va4XrRuxuPka2zDIIzkCF/B3tzK19ydEgvDZ3etiKHSj73FcPbMo/0JOv
bIcB9aCAtMz8Kbde5LOQKmQl/iQp+7KnpVbZOyb4Vx7dYJ+M+mbVCWZAG7aHiwHxQv/zwvzjhoYz
4hXq7wGusEN/3JYAQLvcpzEaSiAQ4wDzCDoXJYTLNoklQglp3u8gEWgh2/Cnkj6u61uLzyQNCW8y
nr4S2YZXbCkQ2PDgUsm4wFxndyj/+jG2Uskia2ZXgxVQpYtAj8K/ty/3fLORcbWkkNsPvEkWJr/W
vv1yOKTUpwcEvhqhMpIp3mRAv+nYhc7AyzxVKPbVSbLpuYEpdsgQDNFNrsDGF5RQO9nDBVqmtx0M
dbzuRkl4Pl/XTzg/dsHTXj9T/XoiK4HCw5xc3mzVGZw+seJKdzoYgtbT4DCjdNYlZ4kwL2Nb8lRK
eoIriDTTcLIylY7YuhbhXEcX0JJeJRhEscY2teJ/UMrSOMtznqHwjnFqj1tNY1rDS8iyFmRnzcCl
qE4EedgHjDsVLeY4PbcvtF3Ewj5chTVVvxP+jusfT9kmWzGSBfb86tvQth4eVOx9O54Db+su29xI
ZZQ65Ajwr+9lzfGdswyevR6r1iiR2c4r//LltEAoS1QwOZ5f7AMQ4qllT9qEvLwYMnx9gbjVCydK
csjvfVxzQEs6CiCHg3CtMrSri9EV0Wu/Ai+rL1j/dj+raoJVWKaR2+KfeB5duF7oPwWIrotT3jd7
yyIB+Na6xGOXVX9cVloKiDnjZEspR5nUlU86V4Nu3HhcFx/d89h3BDLTMctPeg1b8wvQNsSzb7KH
E78+h/xIyr8WMuElVeq5HnZLVbr851dMQ/IK4jRzx5y8MhmIdlSB/A+jKRMyWszhkkB8gR+hpB7b
BOb8e4z2msf6QdS90y4xf3f/AIhXHDQIr3IwcnZIFsiFJiLKJ62vbcT/0lzh24034OPG/wsN9fc8
MCG1vAm3fCGZESTuW6OscXY6E1TzwmIpputONIPCzHiTqt1H1Y5Xq8FzOME9L1NttRDhters2yEB
kxu3blD/N+g8nUh3+fxH7mrlWVlkHjxiGfb8C5OdmLMQI8HmXimeGUEAApVHDt8TaGshNOOzUYdo
lJkYIaO9MC0ELKryWl8xsh/rkmNfCuaZssKkwBCMGrKlqaE8vVqvYp1+hx9WMKQ7T1u/3gyooZQT
wl7hoQFyi/6i8bArfzALeHvocxfKNn1WVdLJXZLzI8HIytT9UrS+rS2S/sditRSs37r2V7FQkOnw
vsGbzxYbFQLnD73OpO8/pb+ckHUQVHqFAAQ0arQcYBySaxkAk5q2IxMIA8Wpb51nWrEvIZq9dNrr
ZmGJIByUUnaAjIFnpoIThZPv4Eie5y2BAfBYc09Z4xgOWGnL4m1LDNKYVf3+B+sa4t/1IVdeC8Ro
ozO7IJDAM11c5dgw43dy45NOtn3hzi2wvP+cApQqtZkaPHz/wGaoxCAoKDMoWlP70UKLPNbAYOJC
q2zBhQZ38C1zjWUF2IeZZj5bJYDw8MeslnwR+aXz4/UHKMZEyk4QBpr8oPNpzUkABy9sTAMIgZll
SOX9atrOYZ/CKMQCq+zWhjMlIRtJQOBBpONJO8/yZtaeTHhYQ1zGTOYsJvFuHxzMLqhpw/uJr2O4
C1PcNFftWuQHgrTzTrymN0Uvt8L/NiPNn08vstR87ICeQNm3V/OSDTefjD78MwW8VgFJE5+k8xyG
bhZkgf8Ru8MsC0GEEWE1TG0AXSN7mixo7r9lyAb7cl/RMcspsHQWf5RIf7D4e6HGZ8+s01LIA2hY
NshvQEhFUyXdRnHnT1TebZl5TKroGGs0qPKD3jUh77etise/o7nsOTegViBADXbXcwoc5RB6ypIJ
A4wU3bLgaGqAtca+PLjhJI0wT07dP24/XismDaQlHe72QpqgPxNPzAh08+DpyrjVh+l+NOJsiBP9
yrABMzZqgHMUO3VduPXvOyyubyDOtU46IUi46BcLlqWwfh/AI8Kw//meOEuVUGobPnMRCQ8H/VT/
0T+lvDl+bxrS78vIcvHBaO8Gb0G7e3MO4ZudOiApIxayzPeM6EOxf+PcRFksaQmirJ48kMGmq5ZQ
5lqywcsGBqJCrSES1AFVn+YakWQhpQlbYw8CYhrVu1uSbXzbrGZ0hEcD5cQmISF65LZLjmkRR+w+
sAlMdgte96VfAu+1iOWQ54Z4ag8iw5gOWv5tFbtaGkENJHsrhD2dUpFykM5VBtajXLCU/HTiLmbF
L66WkHMVru/ClbNxcTQSjs2qRPeuuUtWpTG2e7+MxhRw6al46q/dDtfkiGXbUCmeFLUXUjBoBASs
3l6J1p0AtJuEtcj8jO1P+mUoeGikYQHrL7mSu0v+Lu9JKE8oq1MvWzamjV4cG8M4BCUEDKiPpWEa
5UvqVQksXA4gFbmkYBEZLMtgi68RFmuIo2PxCIpdpHpxNXzpE08NGSKYrjK7Y6PoWPgin8YgT1bZ
ViJ3t//1EPLv9KFmvQmkHn73ZYahETyJD5pbkd7QdhEcN7Bjp4BPDowpTioAoRmhALTBdzTdeP0/
+ln9h57zjo83g6WF1jaUsywE6lzA28FN5/lJ8tUFul/tWcEAs+ZiiHsv7hbHpoaSKigo0LJGDR18
0EHP05GDgwdulpMbmbsTneQMaBwZk+/oTwFi8jPwSRQQNKj2PJhDlTmiXWEe33Sa/NP6oa0MiVcu
wZp0UcEdznLXuDcOX9S+cyIIkojoy+RkJE+j04Oqq1jYUhQznxy1nDAunr8un6WDGokUnioLovYA
yq1VmPtxjMvTtNyDhtWXJjrtPwVv/lGaw1JENdczaWYVDFjpN7Jb8yFGEctEIfm3uIh7aKkc8XBr
HD8hCJRp0YF44G9atqPEeatpJk8OT/PCzaxlUbj5OJxVoByYWeJZpyMIY7DMerunT8Co4avgWKqp
DOexgEbRLsFJIHoVR1geZZtrJP6LA0vNF+I+bcVZnkW+GeXZ7k8UZ3XhPQ+BkNdgIfm8yRtgzQl8
oqfiurrCWJhcY/yq+FiUbAyTdHx5yj11yeexYbWX0gT6Ct5jBbdnfS00dXOOnxoh6kQhrW7n/nXl
NobzEITiuUQTGdZkFlCZP6z5sX7FWs7noZ9hUm+SmwyBd6SzA6JJ2B1SeFuO7RjEp4FMuxn9yQZQ
qZVlpizOWJ21TWoYbVqYa4nvVD6nqg4G1ARHpM4ebDD2la0bTIgwqmeZghDGRo0zeHVs5YDmVFdO
VpwLoU0mMPynF6MdSH4LsfY4oSbi4JmHC/d5C/KC3hC9HPD55JzKaoq6/OvbkVYTeTl/QHEiZNsM
kQLx2qmDE4pZkSy5I0xImFO2zEDdU5Ayuim6mzyN9KoxqPRakdK9XA7ZFVDJvobL4shfQrV0i4SB
ihjlYo+DEQATv2owUhAbbDM+7LQpb37O+olQpXZtCuoPX9lfQp2O+GBflDKaIU0iCRTkzh19gHqW
Fndgcp0aJ+3tIoaheTIZx3DeVzWmR1HQUc3Q8VJW5HJnpJ0AtOZuE77FIbIx2jVa7nHh8BZEbCnK
Yend6kJfrmkSpULdveRNEtv+LC77USmtkCmeaRFn6PPziV3AOpmepi+zDrpam9Dc1PrRbHP7hFXp
0GjieIWdIVR0W0gOuhn0MHQHI+EultqyD4Y0wU/IqJEXsqQC0IXNisNaFUug4tKE9bg20OOGsn4j
4gWs8ma1KwxgvD+/b5IG8CJ9t0d2t8B9vf+XPq1y41D19eVA/ztc8ZHBp2jySU8LZeC1nN6gbYLK
wg6c5MFhMXsG87vn3bcs/fWUfTqcN33YqhhmnILmDDNq7Z+nTAjDZQrQJ2ZTpMh2HdNxQBGOC2oQ
vEL26LkazJFyvgqo5lCfn3pE08lDafe1uQ2AenrydbEpzPOzx7ocgz4d4/9LHxFD7tUuWmQXp5wX
aCYLNQ5rLpslDHpUe5SbpX4vcLt1icT6AbhtEc5zv3urYjwPLQchZZOZyc+UBzSBYsmV0hAhECAi
R0GEeaedAYsd5T2H98vd0Fg/T6QM00O014WEhr6SsH6TPTo83g0NbLpDLBVmSmU1SoN0XeRUB58W
qIzF7cl+nBLa2zW4Y3HufgbUYLsICDl8VS+stshRRfJMvH/hCHN2TLi9ULvB2U1yqXTJEPGQNP4R
9sCknB8pi+XQn99jmEJD4RGfCXFoMrpgpYlB89ip59hAceDWat0Lm1iDZIx9bm0UDkpZKc9Jm5ZT
/nVRZ8iUi4oQ1rgzx9uzZDFZkvO8Q/Bg8h1FJxnu1yKOmlzNEkdyeRtsOu0URgKrt4n55Te5JwIP
mK+T5/zZ/xuiiaVZi3XfkCzirbPWWqdp2oRGsiMjpIdsE0BD/bu2fh3115yGMsxt/1NnXtpqRkeN
lfuFdaTVCg0Z8SPxXjycdnjXUGyKtuZ3uqYWoBeTDJy8rWBPQHQo369zd8XAcKYmL5XhGkjgUM/n
yS0JPLsVS0bd/TFSS4jxRxK0aiX4Kb0VFHBx5Fzz9xf12deStZhV/9VZbjiBacVsF4ew3URxO2lG
ryaYczW/GxVWufN7oxfo8C60NiApOSgi+Fuk61PgDJ+x0iEHNA2yM0moa1P2hLAXQFxweu02hSbo
1FX5qyQVmGJuxMos48/3d9xX1ZXbr/oeZSCdZHsNU0R0Ws+WH+uM3mbxiD9wDd3TDSJU9W/LvQfy
itxrqlYt9PxMfSJvunLNa7QNLmXFIvXf5lPTXntrNoXH3fQ5uwtUt5fSxnYVthEB55CPYclGUU31
25tGHxqr1IljekyvLp/oQnKfQbvkcDgy2XZq/h6e/w7i5nagR3qDNai6K6dPr95T40fFzcnwQ/zB
dwsNZez2MmDzeIvhsZrlmWwY4AuTiSA4Ss/2bA9Nit1UyL+EvHMajpuaJFyzB2XbiATj+cHbGSBo
UyBdbTAwf7hApu2DOx1q/bl/Hc822VEvXAeQr4ZDUcOY3LElabd1/eC7HSuE3TbDasZfIbVLDTNX
47lFGbrQJYpmZVg7Sr+DMBCb0e4Aa+NctUyA1V16wy1vf+cDIISyfFQe6NboStLVxZo6K7hJA+Mk
ckyJPJDxpC2eBiWTIKMGXGIhQNWYZvpX0vhVxzFYDA6X4kzYUC6l8aUBWcaZgWG157lBeAENoUF1
6rjV/1/RFyAMSySdt67W+NU0OVyIUE013iA5xgcdigYqTskomrEy29zIO2SsLsfVmHFGDHzDOfdK
JhzDz6bTvRg0vHpZ3E1/CN0FSFoBod9RInS9VrX44Wi+ald3gGPtthM5WUaL4b4C5PRkfOfLUpht
8O+yKigvFE7FV0VPrRPYqtroAOoU+W4x9tE0qC254o8FgHfMX3TXSNE3sUVHBhU2A4yx5LZt1HMf
7ZVXS8dHwx1KtsPZTryqBNIUXyPfH5Utg03oTDxDCDSLZQywtyBhoCil0VZxHgkXnO+WEPfx6Wvv
CpSAqLxtkIO1IGwOkEhMhBUyWUsOTgyuQkfAWUW4kx+6aDx3jdfS5EDbbUVDMxfFi84qroyOK33p
ccyQSzLDr7uGPvVpwWAqdQjPMKIvShxZJ3zU9LIIjA+tATrtDbSPtUD0LcHx6zAz9HeZFYpgLlvy
+1l1DiX7QDrNBLZEuZfIrtaNDZb1hZ2S+RnHnl1VhlG5lIUoLmW6MuVXNsglPWeev0gPQPnwrkZX
hSbq3aDhEpNAe040DCYNuBWV//cBTftaup3/ymmEiATU91OE4hqoBqFxiCfQdVpSJqPthjon5wHj
+iHbL5Hk2mhqahMe0PhTMWJ1wboJ7d++CR/GNP1iopu7akviizuykx8oFWwUjA7Ky/0csrt9yjql
GQoUL5AkivLQa6hlqeEmArq3Lo7FykVmKhGT0PehnoH7J+D+alI98qvj7CVD3gn2eJ4ur+7qJdOV
dHe45cwMn8r5JK5IAxbwGwXKMZn+lC3emsbSYi7AsYMSGCBf7ORQofOHsKd5EZ1HMYVKmOuQtnqk
0pP7YRDNobs1epWd8IrlxUWcNqjsL8VcOH6xbHkYOS8GrNecQ0S9Kam1UDVelVFCuCtBgCGaNBQk
T8lp78eEhI7L92UF3Qv8ZbtjnCJsDSuX0jWqXQCvMGsuUkPxzmfYkqADcHbYpB6DYS401vmlZ0DO
SWxL7lj/6rg4uxI+cXMvUjGFsS0OUUKSZ3/XGyCLNXUN2DpqkcskarwY+2y9QYbWhpLKjJEpQTJw
bqSzLeKYQttoACxCBOWsJ2bvsRDMue753nZp1R+xvOwUfXpwffj3sQncDGDbulGSwsVzCUTUHV01
FQIxdin+wzozUQXb1dOqSDXxD6vDfRr5nvC3XCEFWeew0aOTEKD/Gww9BeMLyGS+yUhQdy+eSa8d
fjhZI8cYq5gCgtkqSTz6z/6Af+q5XGhUlP9cks0rX1A5o911zbagvPC/Uzj8fQq/P3bGU3G6zvi5
4IWZT4uC+sKq5rNY5+8EJbyyMl/W0aUlDfsd9UHwjsraRu5K+VXg2deaxPtaXsQ5Copewt1Wwp/G
vzzrtkuu7d5CDsLNtCCMztdez1lX10wMgYQ0J+h1RHOS8LulO1BFwenee1OCahAJM2j47cfAZaqe
1tjpLgNN/t6MT2y0OlgN9OaJXm8Hu8w9KQahOcSvJZHVxq7pYsFO9Yd/s5cCABCbZX7at3xkYgeT
g8aqJccM62VadQ1IsjeQiYQpVKKzvYMpWT+gfy/cYeEL0ZeVZsb0VFxwkfMjjAXsAxpgrEwzY7l3
mcFYalqOFFBTQy51wgfvXSei2nY0+ergObVAO8YK4k/Yp7YTwGq1GogLnNsfGP0Du4i1NKhNtHX5
Al8WfQxE81+JpJRthLYVJYWqQRfx2TVtPHdq35lg3s/z0ClGzE+h2pFvQAZtzCkF7O3psA4l0Lkr
aNzh2Kq+O+2qhi3kszXk88MdWDirwS42Um1w4Mbg1mL5/S7nJ8A7UCWAjd/GeOUs9by2/6CCZeJ1
KU+VARmtgEdwp8lP9ShhDObQ+isnuFr5Ish07HTO1U+Deq5tZ2FMH/E/z8KjtqvWPM5GbpvXaU2/
XhWoxUspsq/5D6QPbQdYbWdkYu7pY5CzhJ/rT5TsnsDu4Ina3uOwhNLch1yVE1vEbbRb7HYrV4lZ
kK02HWo++Ir4m0lTp+PW5JcIPRRbeaUarBrHMi06Ik/ucNeivERfWwWM+617asvGZ+IpdH/QjIyE
931Sb7IYkmhsVWhb/PAyo09y8P+WPSNZy5smAaDP7xOGmzhU+Ri1jFovKHvJgLgnqE3Z7Maxt2zA
J0sdMpl0dPOsKjAQfJ2p22xntgA2Z3VMUpsRzNRMPD00PoRDDZ86pJ0Vp6BW/fZ8u2ObZfeErvR1
OUuRQIN7KZwiEOgsrZabxHA7gKynIRlsMhlqFUmLmb/ZzFh5KO8uyscfMYT8P3G1llXMAbMt+fzZ
7jyicvD9k86JQu91MBPYTbCDMaisQV4j9Zcd4S5Ub8Cm6XKGni+dk1T1na/HIBQ9CbnfCQmsMOl+
TH6n8sfjmDOOalweDTBkppn4cYTNn13wbSBgYGXMG1SFSZLv2+U/5l/EXyxEbm1c8/wrtm7pAoVA
TrXU14u0N8WpIIEMXHIIvpZzoOrGNnBBJiNznLaIim/zKKI1XuZGZJAk0b/8M0gEnMlcarOKZEHO
O/kFAoPpsGTS2aLEaacGX+pW/v9aFk1D/msUmh8sQNnYhged4zMEJZicC3blxMiWr/aVT8nsLExh
mA7qGRoykfyW+fozUJD0XQUK14y3B5xEozjf+dAuPtrlIy0DJrfbY5a7lLkBLhhSQ4UsU/5vA2m5
jD4QkpGpVUB/5D2ItKJQHUnqdZ0uDiUpXkC/NqSSDo1jqYigQomeqOTcWtk34kUCPOtNPf46SePj
g6dupDtCWc5rw1gCSFckcBBzlD8+5Qe7/Ac7IFIHn+ZSIbG1acUBs58Gp/1ajqgFP/3bIC62kxdx
zLwjzwAGJFElndD28Fb+1+C1vKz6I5zJGNWpEBkV7h9Kx5H1PzxplBYMJ8BFmpD3SXmU55RN7YRb
bu6mYdcU5vSxIFCPPJNfkR66GMuuYrVnDG3KG2oVZdVdZG+l6eKmqxYvLjj4c2Sn/cA3dAaRfer0
9ScGfycGoM9uZ3+JOz6TY0eQoaIfsGAVJBq7GtqceuYQx1mGhSad7Hrm+rE1i9YrQIt6zuQLmBBQ
LG1reF0bXqkxUikJzRVVoGroJ1Syxq4Ab1paEYW+YSEJNZC9+gC6e2uBAtoFPNITd5Wwn9jevYie
sS+ZNQzxdjmKnLtuwLJccnS6EFtzo17NT/+mXCjwL935ClJDrOv/ilXplU83YOilZIVF0SLe0rfs
uMbZk2VnmgOweVPWruwR59YiCiHToDHGdwhFSHi7pUDGE1J1PtdCbrCHcxZ4H5zycV0Bb1PmYD68
s74o/qFbLYIH8s68RxIa1Ub3ohfzzrJ5Ho2RFgTLZS98SKIbDUYi6MhwQpUMfK8lMmHjqt+v25BJ
obGS8m+ZSvNzZHvfe2UrGPttQFIk16xB6yKBbkhXctyc7gvYl7ZzBft2HgmLXklCD/j1VY+Hiijb
bAnLEskfyz0SG0MW9qjw+7bNbda5hyGqAm0tKLxPLEFIr5m7J7dKva5ZMQfalxZk+tPRacZJSgSu
GRZ3JjC8OxFYm5D4Alhc5Xxr9pyqVZ4F51n27TIBaidtxnvH/rKTjiDZEV67dIH0gx5CbQ+/e6uw
JyqNyIoxyH8RUZ5CaHLGyW/Cjmn1YJV4QPPBlV0lwYkzHCwzdaJBSwBPRRwmSmbUwghUuowJir+p
zrx5CYurqI8n1Y2xHRntSSRPzmhYKBXlIyynquUCTP9MrOjVNaQN0sVYbutm2zmRfHl4FDfhXYek
qvZUUflyJ7mVoDtPeVjuQCzT1QqRCAu21chIBz5rgcqEklDegbsRQnP1IAMDOuD81KyY7oDU12x/
n3uEZBoPBDoTmKwXOMHZcaRlART49kBprQCTf72oY47qu56yeHRnxSyPcZon9No5XZPTgxnytjYi
NU0F8Id+3FUBHJbn09PNw7CljI6bqaUQReOtdm25xnILW35iH1QDOpWoz5Ht7Gexped5D/v3YBhs
Ck7yZc0mmEPS8GbFoO7O6nZgKfHjE9xDA70NhWuMX4+/Fr0pLnZuuv7EF8Ba/qaLaxjTSn0WnCfs
A48EX+1oN9WLWYQ4Mfj62fte4Y21mxFwumFNRT8Y2IYQ2ch6a9kXsz2wYoiPzRzSPiT2MxMIcMj2
+W+Gp1fMvc0gZJoNelaocIsuI3QbRuTVt32vh2FKaXHAcGAgskLGTzz5GVOVqm3RiCEE8H8dMXDf
tmckPpyQS2EWMUTYBJr1KwSp3ugdfn8ug2Yy/zEcQDmxIb2WWcTgfhPGy/oMRwxRuF18ZBtx8xPn
I9+Ng+Fin2CLZ9sH+vLUIhL0eUBoXAEW9dFWx28RJmKvej/yY+7Pi69bQa3U0b1Q6ra27/6+eWpF
Fb93m8Mi4bFEw+dAPBmGQS3PPNivzlTido8EsglIGzlHbz9KNeQwu+LR2JsB375P4IqoRrdW8z+4
Wno6fxFfmPYPvzVgs4unMU4k6PtNFhWAaHmMP0f8MPHYp8A6Ls8rSlYsctDM644qshZhVnSVuBDD
6ZmUwl7xckhEmD8jyR1/Zsw8EgQP+iLPIsQHuP7zT63gTIQxlGo9iOlOVc0HfRR0+kMUQuskADKP
YgV8Eec7E8RVlyRD5Rv5RShmeFQydWs1Wq+BDJM2T26ijnTL3bUeJIOsiakvKeQlgv+wCI4NabL7
8WGaqSlClBnUaGvbMlqN0/525JMZ6lnnDgu577uxe1D9BFrdywK0JreOLIZORPU69AFn/N9M+whr
KxNtm0/arMyNVRe2EZV5fyiPY5/H4d6tBI6+68hNZFFinmCOHsXQJruFiLSY2QLbmGYIC5VyekG5
JDIuW2dvEeW6tM1uc8lrr/CkxTV1AVtw4yqvQjpQOsROKDw9hwKcftcs4WXOehVdeROrlS/rHajc
+sckbgIxhnfeu/hj1lHH76bo/qHgZ3+cRIeqX1eZKqenT1Xbztd/DrlO8PrHOKO6UnQKCX6OuErB
AjXs43inVOCkEiCscFsuaXorDKQjUUv/eisfiWj5Rrgjvy7z8XuDZ3JiXxiuJIp5LTGfeLnkuPno
i7inNg02s+M9YNTOR+clvpEQpgAoaOXTEG+yzApybVaLGS2X6xgr7l2eQ3IvpWXgTLn9IOjfVN87
FZoARDTHJSe0me9jIPvTDcQ22Xj3hfnn6fbquwxsJEkD6IvhB6LM34H7vNHjxDRjvGpj5yFaXlW4
B6DYjGkg7BvSy3dIR9Hqffz2+E5VI4RE4flTDkm4+iczvJbvfTm2Qr30KAvftPuM5w4My7+YS06x
eOoCHwaCdQHtlvwsbWWF0qVYyrhXm4dS3Oo21AMx9YtuEXYV5tQG4pjTMQYIvjbTEv3LJL+yT0TN
EG+dLrtCDqCPsQwAUTsMe8IWV9+LAGPsHKnfbrImRSM6yNzMbZ6tHgsJXZOHJtyoapltr5inWv1M
IPr6BDE7WGb0yHbOzkGNGYDPBFu4pd+UfAXwbfv6n7AzZ6mnQxas0GLjeaWIh0F9n2MmiFCUnTvl
coV6TtGywyvJrMfmAFm5i/kheNqo5FNIJu2X1GQooDxweyuEtOCDtP81OJjVm/lxH9nLrSgOaxLR
ibv9bMv1dEFV5xkKdIa3uDACz0jr6eRKqDEaZSzJq5kK+8uQojIVzKfvAiU97miHv9WNfWoLdTg0
xJ4hdFnnAtNNxsM/VLqmm4m7XopVB0bSJmBpER62GYaMkSYqkvrjCDLYrGz/OQfQoBMhbFf6RJX0
U44rUKw615Y8yqKeXRCb4184rCZOMQbmSZ915meg7V0A1ZEJ7WZ7rw9qpPfnx8Z08jPp1T1skXcL
U0BlCNtg5pcDPCff5AkppwhHKPNNVfeY1TFdHQEE64nKvVf7hd2pJm/+lBpb8j58SkgQmpOSdIuC
cBxTOLfLlnse5WRSuRXmoJLpytWObY4gx44mdUEx/yyj9IgLaYJ8qfDV961uzBreBq9agJfSNswa
vMvSKqmoQZfeHnqJMAs/araTYtE0ABZWprUkKew0aHt/x1NI3EXMEm8wcm4eOMv/KJbcSrHmypKB
kYWSfcYzOICob1BjFZqlzLG6kv+pd9g4Yy82b+Q7Mu1GU+zP+fjKaxIME8BnzkjqwtxCDPZuY8k9
jExIq3F1KKSVQKFfq3WrYNRnXtSifnuP7paXfptzNqVQg0RNIE/YhO/uRPLrhINsOIWhqr9CSf31
/AzWv/Nysr9W0FV6EkZvdTG7JreF+Ji6eD+m1Y2OJKR0Ck7f6Ng9qDZO4jCz2VPRACrBm7fCkHyp
GSUJUlWa8YUGn9jAiUrSPxTwnxKlM7wQtKf6y+xEML9K7ZcxtbxGScwAUOty37CWupcldBVmDT2m
K3sburXoc66CA3Av/oNApWyMAZpdR/xPW4rbBQ9dypuyt0coBJBmawjpW1/BVHij3J+io7aQ+3OC
w9OJHLAAp/XjwbSh+pPOhwHXU0uEGkwlTFlc0WrABtnlwThC8Jd/+2FmxYMnXvm9akFPHaZ/IlbU
JyFyNVmDtu8/ClPmvUvmIa8h3pge+g+fb/hnXBuJSqKuhpzLVJhHDAOzWnD1izSclWmHm7wtHM4k
LxyfMHLmP815ZW7J86y0kES5YsuEsI2OZLv6wAp3jTZLmG9HT7vgC/CxGoljigJM8nAEHnUKSmaZ
0OUCCO9/yJ8+C4fFnfPb2EJDqsHBW5vOQhUeKB+bPSexC95H1SxXcLO3jKNZ0liNXArRvWxal1oL
oEyqHxY/ODzIvIifUpI8P+p5M5Lbx+VOgmWJT26lpmvlSddcLb4PTJwYT1i39bGOjWlatoHvV2DW
RVC+pUGIwa5wPDZOopLjWwupak77mjzWxPdfERtEsnymZfIdg2rQEBX/TfdNmmSa2NWqXO1NUGk0
aMNzGBhtS6Xq09+6NYmNU7vIWdjljytTbWYEKkXM0IKRRR62dJp2aDZsoStlqZfL9kGbr1wP6bk2
s6cR9b1CnCHZPsBt3wBlQWX7LMVTHp7jBp6kJ7mPlxeCAzwpLy9PmAHQh8SztRXqU6zcMwubdV5m
Uaju03GPtTYBUB/NXDSj/M4wB/VFraB26Id1G5SazGWHHSuHzDbUuk8FD3y7b1m8DRnj+zCxOLxE
DuRD6PX4ieWgucueMyUM7LzvZSsqBsorbsOxWX5fxq9WpfJMk0Mp71Fpm9qRx0oX8mEaEDLqRXC2
je9f/QF5ACNTFCX714JGDIm4RwOkOG8fdBGTqnP4DjdHoNjuiN4bGq7Q6Xibzevk/+WiQGc4DWTt
zBQdWcYbgUvnplNpYAfT8XksPwba2OdiQhZxQ11kP748wWLIZHNCeIfyB/Wv3sualcqyWWcYW3T3
9RrhXGP/bpX0j1jnGBEovh2OM8oFMSXMRrX4qJZXQPE6yRX1lUfAolxWcJ0eiTuKX9Ztag90wjo9
P0d8Zsp3TC5DO2wfaGuMBZ/nY6UZiOn0q5aOr2t2Er6T7ksjy05hFxs10PEF+v04XDGeal/RBLzT
5SGnQWhY4JOfDGhvWpDh5l1Y97EyrU8uNtpqMsxfOY/X+r5DcuHsxotAG3m3DRjZ2aNUYlmZTE0o
i1i6ZslHat9H9e1laeVFMiFoAWRkQvQSnM7YGLZ4sAEwhVLd8jXNpEKiRuaEj3M3k0g1KS7su82S
hefVJBGidkTaQO3ou0W9ug5/gEMXsseeRnRthQrTDJ5aKcisVTmieezHAHvVEiUkgQ1Xmx0+z0Cn
R3icAjGEq2qh6aWFOrEYSJ1tKmc1SZ8ONqHxsL5NzIeFjsDEBvMuU9jTLKcgKm7OFpxi2szZm237
ERDSOpIsHobHDgqHpUBMcV+7cP0Jfr6lK8o6dZYey8P9o8SsY1cSlTfSa7xzAKwxDLjTY8Qx+ASm
i18IVML1fEhjfqGM4jLRJSrudRcK+A65wS97ltNw4ym2D7nDzHoEhg9rQjw7zsp1iyS6V97CRO8d
sYLohtSN4sBj6dS7pyHys7V2THcwhR+3fycyg3abywSI7GQfzZ/W4bD2NYBnVKy+M//232Ie8pC5
UT2pqsH+dZ0KYSRu/Y19jYDkem8uKLNztLYZKEmA6ZuYHd/9q9w39YGfwWdsrLGwFuYriYxeVFJw
xHfIgEY9o8/mU0BgdThY6CIlNINjGmRaGK8y0tWJriOdkQBWctpIOUZAfi3VJ84OXvbS2uHK7u3Q
zpSXkoC+cBLqWjPzptM5oVylYzbTceCbJb7V+rub5A3LelF5ZA9s6YQn8igkArQgxaB/NcQMV1+M
n0cFvveRBwL85RTV+oaD1qMHoCWHb42m2Ml/+QY6D3pfYtKAaFITMiSVdsXqK7rNcEb7G9jaMUEQ
s8gx+A4cU0BFef2/LzBeaCyKDhNOTZTtTQbriCNe+93V/98xlmfsT1Ij//K3ChdDh6D/ZDuECbwp
1mzFzdNSOliwpAUZ2bJthp5NxvdR6nvWvLTvFR709VlnMQ0Sc/vJDulAITGK4TuazwiuSXmF7L14
ededPEi2lmD3j8kCm/q9IfeFsiqgGSTVRqxbNnN11oSjBszWrgnNDJoNK+4Zd7HCqg3fKzqee2Qd
IZU+qWED3CLhAo9R0frraJPsfbEdIaY7EqW3JVEfzoAM+68EhhuDqTcvlXnYyYN4RT7xUuLbpr3C
aNX1sERPcTKWDREaN/TqHu7qsV8/Iah18qNv9x0p+rIZnUC0iW294Wd8o30Sul8w6ROporF/G6Cf
qH2KhM8URycDowkRVIHjzqNszGQ7SuM+nXYAQMuz7VyJ+YZPkF2OYqM1VJ6YSL7uWc9s52O0hYXX
zSURiH1Xh7xx6RGuIKUtXTGNhVyDV2SVEZhuAyCP75mt7kSfuT1zmHXesnaNiVa3GDxkWAx+XLYq
/7Qk8VekUvqk7PAf9sTTDRebp3DWLu4doeNvlES3djCRPWHjdY0VwRssm/PofcHVBhNZ5Bong1mw
oAR1nGiG1BEHtKZomhyPlZIMY9KtRRCLRAgpqbL71Op04APQ7TlgUDsdR+0A9R0cpof5+e+YAWpX
hm++xFLgsui/ti0tpF4qj/XrTpTfq19e85PDgwCe2Q/r1WWsC2BIUmNhuTfmL/h1nnv3m1ilOC3f
eMnbXxdK2FAN7MAK1aOXzLuDIiCpC01wI3N8blUInPsX1kCMCgdI++3nfBhrsl2OekzZ6w2LqL3D
SSVx39F8D39ypNj2f8HMK49zLl2aHja65jW5z22l/aT6RhG7xnoOr7ldIx8GQdMa+apHeYiIfsAV
rd36SehuA/aDTnpqXgtqwPb7TOgZKajXQTX4nD8Pjj0CwxjRAyiSPLSUb8Jygi9m7HjrKdgjy0D/
5Q2VtFsmHUSdtVW9f5dWqXOd5TYZRcmLlNNvFQhgLWcxf0DIKICwW2svcmXK6DXg7/FaBD8yFE2u
DV8EBbtd7qQbKfJWUAr/C1PGzLAkuvY3u9xHYX8LhbqPyYIU16GH85fNl8eMyL944+NJ+ulRvkNc
gwoU8JhoJgwxLv1YKLABE2w7u1cCBfc34jSqz1ofLqNj8wH0DW7xlelkj4AyX+QNrkHCxwEJ3r98
H33BVnEjM9HKBgBeRltB496kJZaAkNMrkBt9MffuSFh6ZHcIa/VA1E2UMeu9YPUMTruKbilddtsW
T3Q0ho64IliNLS4xg5+slHxHyGcFMwBvd74+bp3dUhnA8nplj74uhdgV4YQEulPNMCTn/iJHGDCy
2mK4DEsHFFqgxHshDXbpH/rH7/XPrvDHVifNSI0JKQrpsr1j4GBo5egeolkJKyWfkXtvQDdGMIb8
4qgpd9eGGalncBMvHLuZZOb4XW+YGfYBns/tYvhWH0+oHHkK1s+E3uNxWiraLawJOsGec+kxI2V4
k3kCGRgvnEdsImvcUIucpapf0RL3ur3GWirFSnlffXKMjpmfo1xlrQ28lkdmPZ1jdM4g/+FH74l4
2Ax4JLyWaCPLTYEgPC0gWbhHfSLQPWiU9VxDosNqXF19ATfaFWyFekXB+EX1QCnILiJC/Ocu77FR
YomFTmbYZpq41CsgScpVObIySor6xEpUMk9a7Ku66sYGfiwfpJsVEl39OgYZrrEt2lTjUKO69bCq
+I9Wnimf3Os9CaI9X7T4DllGAk8x2+xtPWi0FaCPjPO7GKz0sld7vL0BS8Yr2tAQzBuGsiMR4A3g
dyNKM7TGq1+d+bwkFIrEobswJ1peGTBabbJEN8CL5Ir42VJoQyl4bWw1aS5rleCrZ8QgxR4B+wWq
DrW/9VfsfNsMQDRfBZGxuiYouATESTT2N8qBBUxm7dMUS/u226GmYcIIYBws2ZRahdSQyVZ1V0Cc
3GaDu4PyOYeYxHzoqUJ7Ovw+nBaQGGia/qwUhF0Qkadyt3RLenaPin3+gW5Ye3lDm0QG9Jvm8yrb
6afrLkhy6tgIuTFOCHjwTGTMcymVzC2Mmj5GUARKCAk7k5HWh2NHAFnXBtWab6/PecOozp2JNiGN
UqrXCUwM7gtf34ldxOX/0X5A5Rhv+OWygrv0CnsVsezLu/38iEz/O7GpH5b2ctDccog28q8ljHKb
tuaAwiunEEyWOyFBruKuep9wgQ2IMrjwNKbsAum7phUQCEGYHO6hQa/OgwWNuh0dni3BWHrEa+/b
8zre0g+WeNtYL02Tx8gfvui2+xQJxTX/8BaXECTzAEg6yatnGx0dVabWnIw9V+oE5UCg1K/h0/cz
WeYHim2yAIGJXmi8RF1ooTXmWzwIm+ZZQ7iXCt9oLoTpeG8/ddyZsKkzYF98mlXaEHnIb/+APE5x
FxH+vuRIkm+v0brGxRgZkkYJekoWM3Rxkhle6bjO5PjXpMEKCJX7imbI2TUFqJdko7UfN+HBDike
On02Vp4hwIHv+yIda3+aLWQ8nkYpbL0/2o+Yhu/bZ8YBdT0F6SayY/2ikAyvhKK9d2o+A1pvR5t1
UqiEQzhUFJckrt1t8yekqoRPHZBf1tHa74FbBs6O6FTkPHqwNOMb3hchgdUPxPTw1+vKYQbgYu5Q
A7Gb6nKBa8TrKh6qoHOUiLEHp5SMn6G5MdYdyz0dufs7OhSRAn43HDxrHCCTTgw541d1f1LDfOm+
GVWlgkZSQHK8Iw/GBmVSHbjnDuDLLDRFdxtvz7H2VZ79g8RDsyfc8VoDZXJZiv8YaYEAmNpjfQ4g
QtIKI9Q+ZIapCoDeVZt6ZXPKb+mW1CzVV3O6lvBW/OidVthQJUIIhHHtVA9duDBQ09YDMcvfggIw
Y2jAN+U5khAxUaIcW8p5eOQjOPvQQhvCs4Ll/TQ5PbKXD00a7w33bx5rNfzihCXpVRdMJkxe5p/O
bRplQ32jJGxFn8w/adFzS6vEGlybpoZkIyv/Fb4mRpVSaeK8kjlt/9HiwCkX/G7H1jWdeQ4DlHoo
NcypKga/TFCy5VEdJCB1rTyjRs6zvo3NFKa6I6tdRVKfRRzzDM9HCrGUx2Ltbe///t6hWSa71+rC
pPyzthFUEvuVagmapnTPFRDd1tP3RvCcFhn3jJCG2j0I7+T7WbMrk0VhqJaYBPv+sZYTBTAdHUqx
Qd6He+Lmwh1vPiB1bOZJ1AvaM3Ey7xnTwpjZSa0GGHNF+Ie02gvNEVTzGYAdWnqJjWzpfOqbx5ka
Imq/s3EnUb6TKTVUXEgRTC56WnfUxMOF0vYHMUOZ1/Zv27rL3bVKNsumV3rNfPA945VUSnz9YEch
ApMoX5aRfiME7NRvRiOfKOvCLcZZdCY58nuB+nWv7seZAxTKy5P4xtgqGqsVpbmjFvMtqa5o3XYU
CbEissntGjEa7BShbv6bafxDv+ZPyyFgjMxme6HslaKqU9eOuhSwAeEZygf+T2TtFoKfKX7Pkbxv
dC0fbrWV6AOzJg3sI3FqoM+viD6ipSI7x3ZOJ9j4SrZrHaeNkaGAP5F+DAv/ueXJmSJJdmhQMs2V
lVqITipCImdtVwNHYuL9DUFmd+xNIDGNQhbWiTuKEfavEV4TxJT7nDQO9qo9BoPOXuoBh3P2nlSE
Cs/aSeKR6iWSVLRI71K4vqxZwJ6xMibnxfA5idGvkoBylVlYbYEWajkzVEQwCBEhrJiKm6vayrUu
etOz5mW+vDNNcfnyi9z7DdDHRXWB2KtilO4N4r7j+UJ2EL2EHTB3Ep/3bxqLS0OVc/UItpctzKx7
MASCw8XBX0k7Pv8suyRrvIc7A0JbvYYBwLwTZFwSI1OM6O6oU+X81cAdnBQANPkYJjjc1W0l7oD5
lTtP1s370FgPWcxAZv50Owgs8NnAxjIzOP3uYC7e6oaYTBv/z6p0ziBxDAFGaQ/HLgUcbfUaAqRv
vV1PsRvSBZ51d7LmeC3gGKkFG7IH6VcdNkOiT/LNJ5YBV1W+KPt2TFN3Y6xr6np0rSzhs1z4hKoP
6V04+jPJDRZcjqQYapSOMPOc+FTHrx3NZutaVy2QhvLxoyevb5ojd5jwyD9gpAjmmqmetjLokt2Y
IiJDAnF62CnrEQzUdHyWhV06rYi1YIvrJxvgpk+4JTffHR/frnYZxS7opYAhvSy1BrnmzBHYb1bS
+jtOWVyhtl17g34ECiktXnBC8C5NaRC1SpPKt2R0ub01K5bBRez46cQHmjRdvXUJx9Ywo96hZJtq
nBkCWhXSPA+FWyAYNs+a59wfkV2nfxBofvyKmZXd0e7OdWBDyQkjdhicz07c45GFJ0DFbWtxyhgP
2rDN/WN70HTU2pOOcAt3VkhheaYkgDWEAysQ6KBlKLddF+wXp+ODcOkmjnxKTxEoWMon0qao1600
GgqTtY8TibZNDF2Zh/MPw5+4EICH/iPTnUW1uOMvtyC/U1b3w+++gK1gkBvMlBoTIf1MqmRC2rUB
EwNAqgUJiSJcLBWpewVq7YuK+F+XyFwapADpDOQcSaJeFAJ279n0ASQ1OgprpfMSV5msz7rlzsoo
AAa54zGmrocaJhZbMVZSlwsiYCZG8MzHXdYOptcwr6c6W5S0kV4/YYxv+Hi2+DJULwxGjNtuPhIM
4eqbtLjqmPupbw1SNnTGHNfytpcQWA3UjWxM8ox3fQ7ID0JGRRi/Pw+bW+yRZ7lI0Jv/wIurvorx
Hz+FGXoVe86xKriP2Maq5K8TPKr4t4sfJbxayKJso8KDCgOSll2bmSHB6Z1LLppBBMzjhuiLKpBP
L63LI2cS9ecSFDEhePm83d79WjjpnNC89h8Xzb7aJdUUGrIEVkJMnwoEX5Zc6z44wQAoIda891Zn
0K0AyBTCsJSX/gBqV1aEAoA+DoE3c2y9lQ/OodHz0TPRVAzK57vwOdx4XheBwgRrMsWLFioXJ0qp
FdmTRDujC7HsZD6XhBP6MU4HGX9eSP8Bpp2zfRQskjMsXyfzzxSRVKCHmpNxkIQ7mZ+Cv9ANtRwR
3IKUJL0PtS7j/rE3KqqFnmcCg0pPbni+wjZn2vb15FTtZBIwMgEklwSpU83caboUsMyVAsh47LGV
p/Cx8Pvb49DAXRNjA1Dx/z54OzUazKojH7wggkMwnEFMA1M8I5E5DoFpwQWbTYxYjZMXBWeylbZl
IxW5cXBtpFeK4IBFxBWE7jz8EgW5kmDV+mYD+ctL6WCweuydDn8iWehXuy/EFn3jn6lh3l3IPumi
YdafaJkFjTJai5DQxuPRmRFbKCHgNukbQyL97EB4VI6ZOB75KDTN7pz3dGbKUda3F/yEEyFAb/ww
fiyMgPYiaGc1rhUJWJCWV42dog/IN1cLkwmFrt7eC0oRhn/UsMC68K0A5gOknMIwDwtS5VAiuH6e
Bu6JlpJ0u72B92fuud4vTNH95Opdrwl5wmAfzgQyy6NKK6ylC2Iaivhjv5LKY4W0QQrmIVan4RLq
ZyUfFTPHZ2oolVcmTWnyiwvYD/EMM3bVDxyFW1/qSPcyT8Ql1paAuqD/RSkQ5AwvR7v0Z70gP2lq
Q8+ddd26+xCn7zeX7pfkxMv/aXhAkUc1eKVg0wGzow/LwnECCiJA9eTwfUKfthqd7jw5IldT5o2d
9cWmo9H/6eC6+WZ8MKnrRqP0CEX2HdXnsZIuKARAiRPJ3HWhQMLGkcMHxRCjvLxhJrYhjP3zx+T2
RNicYoFkQjeeVOSF4XUjp5eLZ2mEuALJRvsRs0hPXPrN2F9Yo+heCpBK289aC0DYAXE5p9rFUtIz
anOBup260okeIcYLagDkZCo8aT92Zcd9YnBsZjXRLDtdmyj6m7XPKNAshVfh+tGiiQBFsOOeaByi
Aka9h3iZvidcOUUGcmq9jEtronEXM6p8qEZmr3UgmOSlJm85QYzywostgGbjKQtIE9XRxpzUVKRa
jeKWt5nvJ3GDkGxuSHXT/VXlMwVPftk0fSLfGFPLOfEb5GsuvnsXDf8ljK8JY8j2KTSzPMGAulp2
L2COVdsOW5eHJg0DZG786tVs6foamBA907eaRZ92lZHHW6Y6M0tUzavib7L70C0f0Ry7qcuORtap
Flr9v/C1XjmRIh93H8dwQ4lT+2q/VgcDrY586G2n+p+CcofDbsQrivZ3hrekBhhKw4fv9WUalDa2
ptpw0Unfi5D53HDU2+VTYpXPIzX3jGeHSHAvWVWWm0+nKOhilbVnOa8MvMuVekWeL/gmPJ1vNy6/
5paaUCxtq4bbZr+3O3z+pkPsV3dszUMNTCRY6s/3zwTp5Rnyq2r6SXzYWCk9u5VMkeb5q6ygEe/Z
pB+Wu7Aojs380gp1RJasuDTjbvB7Y+eoNJhYvVmp2cx9pQvqL59d1OPFSMNWZQnOdnL1YlY6r2CP
MMjaOx1JcAt4kVacjlokUlheNFw3mUUGumINwlqMKwVE2SJ60LIyT0kysYreONfB0Tqy25XvvlJT
GZLDGjyETo/Wbdn4AnxaPw9zyf/yOFYhkFVxsMgzd0wtVPlFsC+DpvJymhb8Fr3povQDYEjzxPth
WWMmqCfkmBTqNLTO7WQU9rMZ8KE03lig9RUGWX+j7RN+IBrduSsGitel756CFMgDJuBN3C3LF8Fg
t2gYTW7MvtwxjJyR8er0JrsZnTFIpg3oCknt2jr36khADhT1l150gZwvhvfgDGPimS1sxGOIW9RM
u2iqQK/YGvbzOPsG3DAB9E2UaopfdvrdIKtY/xlLd5g1BPZaBa/dmg82+ImekrHsoww4fjUq1JH8
Gw05njcPM7g01xJMlYGnFMNSHgVMhbocm2i2ywugFaUd4I8mANlskhSvXacrqNio4vUi8/PxovOY
lX1fFDypdAOy/4SnIrsizMyHdwjKUV4R1ppJtUWG8i2KcjzNlJg44SdUSF3cJ/705HJmbY18efOV
A3rntxw14StjpfLl0VU5PxavUBWw56aGislNQ7ykVj5po5OlbYTvoOrAs+w+R4zYVAx3r+NsjtS7
7kF/Hn1JJbXetYdpw0fgYDnE9TBHEiYg+BAz8kxBqR+SMUd5FLG9kJ6NQiP9Mt8OQ3hdLO9gPijW
+YXw13BzB5WXNZNKWX9HvHQNhgE2CD3UrEbDdeG8mVfibeZ2t1F9bmBrT+U76kZrFyu/thvc9+/Q
7zrABITnk6XJFc+IE28jSHI8eSb38DSqL0TFUkk+96xbnaUko54O7hTA/nvYGAF4v64RrEFnP5Qw
6c86W5v2mR8GC/5h0Pb2zsuGYH73okykxvQN+7E23gwG0HGYcvvqYwT7SS1wrGsjoZpSwjC42II1
8OdIK6MhAvzLpSyQZ9P25bmw5b4//lak8ui4a18yJPa+Fo7jowwCQDe1CBprv1vG9g6ddugpx4Ic
RKMd/UHSEZHpQhtITcZ00cnneeReHjnUz/VobPsNzWOLoHryBOsgMnMpZ+XLzMDi8Rty22Bc2XEP
gX/6PmmpiWaXaF1S90atwSNnTrpnnBOo630UamZ9sNlFPSKvl+uag5HxPSjSYUZCiMK0/g6lH3aS
IxWp8fWNTittn5rOn4Sy7wYXFvlAP8N0j3OPGbk7vWxC32hfE8xN7gSjT4CgjHSeMOfSQCtsxoOb
I+jsCAZZkbti2RRmgv7VDGkXllf7BFOizQy2MTbGPQX/M14dMO3uJMwEMlClLbguVFuseJUcPpJE
tZVhUDgIjRUXILUQ0S5NAeYbKuR89YpZLFrMPNIMOt44LtT7stnXETLPR3wc/1TqgK9Phr4DDj2b
GJOYagmo71Zs9jvq6pD7gH5Fw/6EW2vK6XDyBJRrKd05sPAfvFi9KmTRjHV9O/yxJ/oQ+F6+n5DC
YaBwY4MJiLU8K//+ru20HZX2bf/5EDPQxe9p1wCboiWRGpQr4fFc8FcCAPylruLdHJgrgZ+I+9VI
jeW/r7o6GRQeREWvuEvWiYt9vsq2RlgDsu1RniTmsxr5SZ1MWML4HqJDm0xlilg1obx9DfhCiYpS
8/kKvT6LD8lO3ihXGkzVeL3vjJxzoSKE9fXdlIQk7W1Tw+u7ZZZQMt784xx7chryfg8+iTnOD0X5
Gnet2zjYdf3/2d2+DKUXlDI82MptPtgy8DevQ2bOkxIVWEwhO9Q8ZAxQDd2rfwI/thSYaoukgY4O
Yhf7BcV0brvsBb2evoUs372AI0YK4ghLjtv5UKkuvHUHriqTWx7CV1IZiiJvIh5r+QKF2j1lRwPx
4PuStdLJ19LozZsf3GjfUJp0nsDPItfse0LnseonIpIjTsr9vqCzf0vqpCw8D1tmsQfWK41ulkI8
k4pIz5hXyjRrR8pfY5cLTWQOR/+VPOerPTPSCF9rAMaYudp61lU9+5RYKqNPQ1evL4q47DVJBJKF
uGMfAmMSPT7xxHpw1AaJxlNm9WXkIAIYm9+rdqPDvHvMq9H4nv9mC5hg4QLm7hlYFprS60qJVUli
GDdaPmdzhDhB3pm66CQNRt6r6LfsjNigYxATCzVasgty5KrS31oj0tYQXz00+s2T2EUy/isqS6H8
hd4araFk1I/AEP9lRQuofMs1kBg1gV3EvIgn4nMV06otr5DwfuiYNDIakd8nbXIGdaha0xDtjUCN
GLEQhBLjtqzfPQ5mtt8F6KKtNVAXcEIUbC3nqjUfVyL7AKbR4tZxSW/YMIVoh75PRsbgjOrJmSjm
tAWs0vtTpAssD+r9MZp9Ec3u+3UkHH18WTsyJkX0N1tGu5rXeV/VckaoDzZ1/KEQu3EO4QHxqwB9
tSbksrECe4BviVj7nrmLcIYLNu2bAZUHPUIqsUehYlmbilq4s81R9CfdYVx78apWG1CzTyNKt+e6
HRE0Hsh5qMIkNdQe7lkYEs/6IntTQK81113XhsI/88kIrQR8vkmZ2UU4HpvPlLxJ2ttRGlr/oA0V
4ospPjlaQT3epWOTX63waTnWcIvMftY+h/Xw0CykxPMV6COiiZkT24cGRWGe2cU8kEwiNkx3d/5+
S9bth8Ui8yRm/4Ovx/w3MclYzyXpls3Ocl0XxgP2xI/Gkpt2ZXG3/S70Du8GVSqWNIx8iRUW32F5
Kbcv+Z+zp39LtoRFJL3UyDIwPhbbZ1LGVNYju3bEQw88zrcc0gOKgIwqcqd0VS65uT/sg/yjT9LL
ECpMPG0RR/h3fs78Ep4PXVL5/xWnVh7lDHmKIj8Mydlm2pT7oLpL9gKe5dD7bBC3K65MgX4DOPYx
UTVk5NWZwGUGYWNa74s96ziDwpCYiORYIy3T8VlS1v4fA5jvjgWenTYBqEdHK7wV7YuX0zg9XLmB
HFXqc4i8C4n3k6Nz2FB1feYgdfpSdeR4eCCHg1JAyR0h+LLIplM31K2WHaV6fUop2xyvI2x0xR45
OOnT9qavH/li7RqIWhLNHwFv+x6f0iS8FMctSA1Lc4ooM8Hn9cmoYdtsoJIRBO1FF5DkNeLM4R6d
CgHMBjYTw6Nu7iGqV9Z78yUzumYeAC7rx8uVpeRrML0guPZmDv5OQ5AFHbXMYiNltL19ZWMxvwBG
qpd5OthiIg5TXXpOHPBEJpW0N5kfe5+KClWuBdUafhfUtcDi3mWPB2s13dmskiV7jy4cvaOSX6mR
oftgyXZD7EE85vepOZWvggvDadXNEbY/QJ29JKJVw6yfRZVYEPaTeABKQluHavsfyP3OAMMzvfSr
UeoRDdFG5i9JXG9WjNJ6tYozbdwcTlt9k3TKjuj4v58hDs0xSXe0GkgcDiu6tIOipiwLLmdgBkdU
uT3BTUFTDH+ZmG3AP00p68mKrTTiOoxKErGkPp299E+Ss7ChvBo2cNDtnb6I6Xod2j3/hpKVCRKt
4k0QZSFIQRYr2nhcayMNzqnR8OifAOZcYG7DJmUIZPNvOBbNKL4E+bZ/npj8fBxYAAhlJNha8yae
aM2NNyt/T4X2FAhA82+KGShJuvV8YfjaiLP0eDwYnhkrV7OnOVilE7l4Y+cIIzCkHpyR0v5LGvgQ
2Ih25Hs0P3opu4sDlvJRwWHtbRd6xnc+NtnAV9QUxc4mBTH44fQVucjUsMrs18Cs+LyNu2mNcxOI
gk/2sdcHjT6gh2YmWYhlyJfKz8XFQrisQdtecbzJs8SW2HgYJj54K16RV+mrl+op4t7/jCryF2oF
k3Zkw9VPd8Aa9UGwO5kr7Tn7SfdHng44FInQxQ/CE8LRYYOaf87ioutzR1Y6W+9JlknT1U8j2m/6
EtpRN8lhGxQYNwJHkVlwh0sqc3fEYuGmXZ9Rg3npwKl8GEgCHzURSe4mTul7fpa3LbGsCg+8EL3x
BFbfo7SJTThL2Vv2VGPUOMWoIU1tSIGvrxtuBw/2m2rcIdfLFoPgxvmZD4UJlrreWUX0o3HtUJ69
a/sw5zM9C0u0T96f5c62ajYaOH2nG3ZP0knYMbzDw+YPx8eWcilLxxmKWpyuX+ysC6llrvVdD26+
7yVxVoLfMANOMQmV6r3gGodzlXImKOMy7lRdw+t5JHLZulITlv8ulFaCrUe092RfKu46eyGvCuVX
MyijEMKHOy/66/+F+3wxaiDrQWwKHCpgXnhLEmiqm2n2xdKjn6dWWUOonVkmdASBUyAUMSB5sttH
svu4xglvNo1OTeN6FL/M0YvtB4aH612Pr98PeGXyPApYYxiGpGAi0ERfuHeO7UNpxQgrSO12ogO0
FzxHgUocEr9eeH2RsYGtf0uIpFGoskvlkLSxpXjcgBY7Uz7NGCXxl1hs06hyeWnwmYCXUcFNDWGe
PXEiuQ4h+07gw9Hti36QJ/1RWnUahVy1evFVPIF87rEmR9jvPTEkUeDXIsTE6mwpP0DwOY54po0o
tr3rIFhh8GKVqJWHsGGjN3OecIvECYQq19vVPhJNrJI90D91b0AoZR5npRk2O2ZUWE8HtQ0FkWk6
g8iasfgQJeKmPUORxzqEADcZklrLMMhlE+FRUmwoAgTTWr22oK8ReePxLumuOcgSwiVsRxtjPl2Y
dSZuxbhRbKXKvtH1u0mUYsXXwO6rk4YtMDSms61YUfFawyKZK4qNRbg5elMnZG2CNaRclIUV6JKg
02QGURLqvBJmpKwv88PHMVDuLlWoUd3bjDb7edG+1KcqjOFXWn4jJ+HpAR4wGoFY1oGkYG4wJXIz
4z7DHLSu/hmXpEbDjZNfapzjVR0LUxitZkq2o/NGrrOj+0Qk3t56WviymDglyrINr9voo20HzTcd
XP0OVimANLtLcIFjS7QT03WTHBZ/6BItjJlQvaXA3lZbBvQbd8PwuMXdw7RL4t6CtEcEm7rG2jxP
FEhnObqJH2ZRwCnibea3Bl+y6WnrAvFk+p+1i3jb2as4sdvYUcSDnPOPNRnKMPmV56RYkPTCx4I+
IJ+a4kGwKA0QmFnoeTDDEQUAXtka4QsLwPjqRylx1d0LckdUrNTNvCfKCBfp88415yvIU4JBxoYy
nQY5WyFpSLU6uBa/GDJJcAmCSyQjsrAYwx3AMkBwUZzrbdWy49UK5aclgvQ/egJ8TSUy1t6QzxtO
glT5sMgaHOHdHdZSyISMqa0CrPZFrwWqFTme2vkWBvOra27YAOsfGbhabWFm2pyyI0hLQ5bUlVwv
V6OxWCSB2UMFa62ZSWaISXp3Vn/yQAtHMEgxnLFBAGPAxYgSuWHaCo3WCp5GfciQ7vUMum81jJU+
2A/C6rJtpt7XPtL+wi3zIVpoTcqmEJpV+TAum3uEVyf+daYv068yVzac1EeqaMuX//YYzSmtLnfM
68ZNNozYpimLKkvwxaANl2TgY8lcexBlUmQ1PqCs5M5xDCrs/mhn05SXo63lPFoiF50LlZ11jdLP
igVI2FHEpwAoC97zKz9WXclJqmEY4AzZo5qEQ3M7ddIKPvw/NVEQqOKRAZm2YCJgxwB68RjFfsGp
8sGW7Y3x6AcPWrmzVElMY+btJjiRg84t9Xw8Zxwpoo/XVrtTP2ia6gwMP0Zr2kGsoP9aaNE1IILG
Ay4sn5oPOufBMyWie0Ua3L4kqTow2h1miyD6tPAFVon43xgUPfbnjkpWiK7PrTxdmNcdNjaPgbkC
kvJZuQG/j51SaBYAezmGWNd6QEFmuVkmOcsqVOMSr+TSsCNfKpVuxq4gFoet7hKyGdpye4K+LBId
mDiK4/o7tYUIU3WodArH8KyTgjnN12trPVSAzQaJX6UmmL/z0siJFzCKlsgyisAex6MJT8Uwl5lo
33l6AYoOGW8UfzudmGZY09UFo+w/D3shE8H1rdJU1SjIDci/T0unrOEqd0ejXnAs/qbXklmXLPGv
YkqB1IZOoX9ZEpQTEniEruEzQ2mFIWri7luqVDP9Gob5j5lx1Wq5TkKP9sduZw8XQuJd59E1rZZb
uZYMbZ3SQi6E/CIBtpsesX7r9Xq09YkOXb/oiFKgdeFVeexUQwHq4glMXU+vkIMRYUecyDRY77OU
/X5QnNTaZzU7/DxDPaKVxY8Ub3V5Y1l6al+9zeXEofWuWTpC793VTmBwp2byK1HwTSJBhkg35n9/
71jUBvsNCQWH1UgVB8SCLi6JTUeyuFQl6Gs+xKEjBXIpewbC/mzE1CNvwYMA6TN9l5Xs6rrlm7vQ
XV3ncguRxAbBHXSBREymtMqNP0/YpOxbIw1ERTkv/pyyfYn+PuAhwxLlAzGpCxxjKdXi5ADS4Z4Q
OE+/M0ll4CVRbCSRuPjAsuarf4Eby8zUCVmixHJvHLt8bPpZYki2Tfv5Utsv9fJDgzaXaHqLlqlT
w3CK1jZZYP7ZY2QwxhNwlygoKvUHHJyAmWARKwDnqjiPnyob8ql6PnN+V/dxtmy+8L4qztnEv0qP
Qdku7m3/XfsaOnb9MoflLRxzLR8F3B07JKtmNkIr40YXt3poc8dYVwc6YMZRKGAowwC5DgXVP44r
pVzrK/7oYX+7rIDmc4FbehpWU0UOsPccbPaLtq4iGn+k/ntinD9YUMLhNPCAHDbpKwOJOyNl4cs5
+mxsIQDIzM27Oc9VljOJZG3WHjyk/+pnXMiUktGe2krP4wBViDUJRnASmGmx3Fm2vrPq/Fl2he/n
ZEUCOM2ZETfwd6qyPaABxWg3+lc3PtVC9A7nimX30jUn2dXv1MJtAO/Zx3Rh+tslg/Z2igtlTZib
1PftjQK6wQNdaFDHBHS5ThLKuB788o8cmPCqX9+xiPty0QEsCS3tuMvSKe35WYb6vj5rwDXTVvp4
SgU17R5aftmEOUhWerGJ/hZenLSsQEgJDQngv1n14N0VSN/XJNJRLlxzVRRQtocYVqPEbIVn8oof
UwXSC5yHhcW2LebMFsQlFTevHUOhTwjHd42CPk0PX7xsFh+sR7NoAguARLixb+1LpMzBP5BZ6NCZ
l2te+VC0k5NpsDHT0Yn/UkjuATnOSw/bpN/m+w8Vaye4ezGQ+MpnnBYdRlIivze48S6IfO8YJPD8
N1P8EAsLpkLHqryGHOsJR2e3Va1pMWvWsjV0bhbVfElJjjbnT818ZxBoGd++X9lODJpFO3iSyqv+
Nlb9OCWzEB8FzufNNjpB8u8WPC3KAkCQ0NpWVsCREBbA248zFJga/8EVQRMpWpmeYm/xXbIm4mtf
juTxr2lVJMIQgm+ZR/78xkN2mAUTzrafzaCYRh64fRBoq8QBP+UKJ5CcjNLKZYuSW+3g6ylVTsOY
v/o/Wn0NMJRpegNPVBHVT95+xDqOXvsFDndn4W1xNW9xhs6OCFgm82UeWcU+J4K3DvRwUrGQtiks
E+P5/XFw4Ecf/QMdpBRPzNcXVfqSVlrNn83vx/tGNvcYcWsyLMY/bih/HbDq8Xx+0HSYNLBwJdya
tf9416Yp2aNkYLeIjU3nsEXGFHqnSaauDfbD/8hYAvHELS/wh92sii57SWgNitg9aDdnsCz4mTnY
4vF681RDllPb8JmZb6sIsmzHW0bQ1dD7XN6EdHrOt4CJ7dIn+AnX1idTAqV3AyyxXi1wcAq217Bt
JclinpDCd2vjjtxaS5bdWfA0S/eA7s8v5K/31NTz8eJfvnM5VTLbIk0uDAMNfxzo8prprF1GICUr
fJXexY5EC+XmwSyYaEpdl0sUlA8utUwRHn7Rl20RjUQlYJ0Tpa3TfybIn6MjxhshY2aYe7PI+s3P
D31oKzcPHRNaKVCyQK1R6k9YHlpqnzxJoAfXLAehgCim+EMTUgsAKV84yR/UrLTsYNV8KKr2TS3K
Auc/HvDpyTNYVPZM+9YejywvU8fEa5kpS1/X5KHGxVka6KqdswC4XuXSB3wqLOKaekDyx/a9DRTT
B38zzRioYoLRpzJ4R0tRUgA+Qg8NnffK2TAh6ZGzKMyuZlT5YuFZPSxx3pcyxOzt8EgDiL4JIBs8
4Lf8TY6Uqm3i+6qgQjU2Z0Uz0N5aMsLKwExOOtWji6Ta0a7P0O7mh2FpZQY8OiNY8V+AIbRZdQ1E
e2qgSxX6DSekSJrdVn+vzRBzZ19mgsyI/r0qWBGJFrKO4PjzuMjjyq7i6PGtEyE/y42phk0KH4Dq
yBQ4J6cO4HjXlBR+6VNxj/sMA0HvjyRSZDX6K+/k5+Atfoe8V7XrKiUXxMfn3BkAzuCSVbVMYJef
KxJEubITzQhCzr3bTHA/AI/joTFnwNgUDQlR0dluShrNACp7mmP/1spLUqYlpifDTd/6ci1D/i6V
RbteqQrJzbumcEx+oh895utaG2lpY2uFR6aw2U8PkrVM+2cTO+m2b7ICga40buWIvNdsD3vUNTXj
TmEdtSMC94EE+B5SvV56wmwGbxJ1+PP3pDTfvCFJYgNLhY/xxzmtDyQmriX64/sFlNEUMPnTZwGo
ts7dVjLIuqhA9jfHXYUZKOoYb+w79eaZYyTYRiPD2zbJf1ilHmrkz267y8dbnHAbbrS3bpWAac69
V8g4a5RDAVVo6pW4OA3FIHrveZmGQGneVs4kgf8PFxwMK3+r6mBI4WD5wT6ke9X30PGUYOtZ8TTT
+Q9dbkztnC7x9ybjaZndorTpLUPK68x3elHqVVkRCSfuT2YQpBs8oVjnqZK8zEFza95AHM7OLO/O
cHYJndckEBa3ZeZOTprqBO4i+aS8KOul9rXF24HPrQPKGGTmgORZmYbGjhAat9kyK28SS9STApbY
0dkJjhOWaHKSU6A/2RSR6OKTQ5so/kNgae1dP9I9rXLcBLfwwPUZ6RS1iARdLZ5g9jFQ7cJNoRpL
gd6wavktosyH07zbWj0rFbO2o//Ny3n9jGdOwY1RRoNtSTFt4dHtXlCgNxr4quMKp6SPW9M2bh0q
fDgt5TU/hcaRZJZwIvZJ7Ot6NXIN399Twd1l3aI8zlK8mmjiaaQrOVFabQKDbDr+t6YoOFxKzd+w
5SMml1Ka0Bb53T0hGYiJNdbFrqhEv3dVqiO5Nm05Gtl8ahfSBO3E3QD0AhFa6N6Cze3VH4nPAq7I
qmT2S7mNWvS1ne3rIJJvEJR2+dqNQnXa7mX0bx6/4KhK3BmXtoCw6MiFQcqVktbhDIdnofrtG2Iz
aXyq6lxOUnko4/bf/GBOcb2QLJOG5DEIJxYYf5MfAQ8cUnXk0zzZb1lonmFuHFEXPOcJ3wvnU/Hr
CAzc1ZGMkAkvcQUbwkOSHgKA/Adej2k7BKCRoZQugP0OJ7H2eqpdJCscpPzYy+DgIDgP3DdxyKvH
xl5KDjwBWFKEqCaBENEzEHDt69JZ1AtmSC98hFRcRHk8CMYD1PGFxvLovXkEf3Zzmt5gO+VXUdRS
N201WSfDx3YUFysjQOI8C4bzRa4uhNzbEtBQuJqcrq1C2yNUo5sw08YcZvl01jMc3PkKEiNmAliE
6IKpDEIxo4KOTWBELMssU7it7SGe1h3i9DcqzbRv9k302JUdaq280Vm02vrQwO3Eo0mIuIiweAcp
k/1nMarmELizPrRYZ6c0K6jfxRgojJTN5f+R0zSpdoTAxLRSNMrmfDzx8KISXo9mSY0WQ/Kh2Ott
jjrYriHeqyAxCl4YrpXeKDx+rsFvmDs+OuHYPl6vcKKYxlQKiEzKhodFS/k88vJexIerzNKwudFl
ZhyqhYnqbWnHWBnNjIN/EekmWJgk4LvLyiu5DF+w/+Pwg3QpvIkZvxss+zngkJfzLYVltHoDXiJj
L5k/9YjbMRNBjd6lJCudNNxdKG7sYT3tnhkY2hNkkR3VhvGjbWJLMytpC0L1UBNmExlJKMv9R3MG
UpqYfvs5hJm7FWKnOrmO+cpvvPmnlHgONBSuZC6uOUmE/g4/4TAiTtOxBZT3MmCd0aq8UOWAwnmb
7LD2+sXRON81abMmxAEELtV6Xh/kk4b/cpiDpxOOLGP+z6swM2Pic+Z8PtrF2Fq9nK+gDeMSFj7b
qUsVGWcYWiHHiWJpZ0SCHNg01u0PqNUMTJZMnERYS65DwALnv2gRat/EZOdKEKqCzEwSsf9FOo6X
ps+POZ8IsKSS1bG6r7HIK/nKtDfemYCcFNsRWhikf5T/9rzTnfsmsc5ncfnzrA5eDPZxvF+Dspbc
h3JVJkQLUxhkTWpZ76GgjNUepou+bOCbRasmG8upDVkvOluyikkAXmmMo+qP1bkSITQVT7yeCHpa
TKoIFtHW2xcDztXmOTjX6FtmTLcaUSsaCa0GzM9NJrtNWTwD15mv7ap5UsAovnnfQW+vB/EH8GL4
1JTGn2clFcOYnjVRrl5ALt55wcs+w81mqJdT3XXZvRCySZSlFJy8p4vOguQF7ukzVGKDf8z4E4Nv
LkJL9fBMu8DQM7ERRafF3taXjJV8vmTX54cG7SyyvCS1V2yY3EaFPbVPAK1Pk3SuPHkn4SO+M4r8
rvXBf7rxx4zy66svc+02SeKBFeSNm/N69FOclG1WpqGp3inSma9TcYwfwXxWD3xYHNn+WvqF0Gl8
qjYl3qZlR8Xs2vu/fX7+a//KKm9KYOgGfTDNH5c+5TfjjpKWkoZ54Pa55w44WVOdFLbb7S8obQeK
g9n+0j9Ms+dcQ+oQudIbqt7NXjmYbIiCg9gzyRhvTK6uAZmagoaR0ZgOWB8LKmDJKk+wUkPYpyQe
JzKJAV7iRHtWj9zGqOXEGN4hg0vi2TrvailZRaeb/xqZjq4isIZ193tQXVFEl5zoS3rZ+fPDlkQ2
v4cxBihwts+OYBfffmaPsK+jV/GGpQm/xr6aFtswwpaFvEJhkp3kedxCGUGzyPdv0W/0DUe42REf
O7xFkOfqWqTZ4Y3rgqO81dMaeI90k5xQecF15JSttoGRzg1hnnlKTHCapAVMICiroo6/bIr8W462
UIaZsYsyoz13c7YIo4jaAp20pSPraZSQtVc+7X2E7047ROLbMEP6PEQcZZcTRqQy+uF2aU/66E64
L4Z7cDDg7Pv3PWVCPXVJ1SF9KEi4EdKS+Lq4dDuXQQeXRQHGwHfk3EwoNfPXhBZiEPe5j7V+BMG9
TBdG0FOY3dJZLwX9l/3j+2QblV9gK98CllcDSj6FC5iGZysdpiRrsvRUDSF6F1wTez8c/RvE89/W
1RKKReYEW84XMjhlrZtdQeiN2z42D851OxWnRt7wLfhKfm4lWs71oKo+dooJQ2V7t8Qx1+6kh3I9
LUjhVXMi88iyl1EiUy0l2Uj7aRYO4ql4iwypZvuXlWxjrlVN/gIA+RX2YrHL2Vs+u+rQ2wDmj8sW
HQMM2koMemqqYeQmyklCPcsbVLyuK19uKEjedmvJt4NqJdyZCubhN1fW9eu55sUQ6VEbZICGWufn
XWDb9UsE3i2Lcx/TMziaJaPO7nnJxOvb213FuM2YJ5Xybc46kcchieVCpgqxfPOY04ohs/Om90Ii
P9agHr+No6v770FkreMvMpUwlx2QsjwalyVh9zJOvcLZtD85bh8S4bfrVvH62hxBYY7a1tkrtYrZ
hitZ5PpoSKT6PXeLGX3Pjdf/5ahuISybXlEmT0dKfr0r47N6KVf1rsINqN+TYq1kGW0Y/GNDIqRm
UEDgibS4trZ3tuTF8QcM58WT4nyYyQUn4aEFbxfkrOjLESoHYOgXqc0I7WH+mlFMVB4fll8/BZUO
Rv5iDHyD1W9116kLQaHsAjpJgWJl5hqHh8Qs56NJgJKu9T+Rv9MPM7yI3DX5G9hluXfXfsN4+QBP
VzgpfClDtyGyVRspY0MlKi+2CZVvndRfnj9y6zq01GgWWAiltPzLXfJ0iybbcruaA417+bVW2HrC
fyWHc8DmbqTDWBA688r5XGiB7BmlqTkxE5zJrLkQD+LnK6psy46XIiEEOAYZRpHt2t82DtRdzbqW
ViRu6fOU7Q9bZXHeby+8ATahtWpyT9s5PGrfT+nhBcT1V0FOPIE6KVTWwBxmVCBTvaeRHCz+d8ns
hMqH8+Ojdf5OW0AaF2j2Oay42LwybTmatMePtl4sHYJECPHjaIltbc77UeP/70FSDbxJhmU38xVF
tJLM0XBakN9M2TffmJaHrr5wnPhIjAu36c+KOvbFd9MSu9qq9rEZl0zaADWQorLZ//4d55I9tntn
iCj768JMtipu9YRIdZdrvnWrtbjV1NgGmOtw9iovMUSRVx5iPr/2atA9Y10dhxepqxqsZKhjnfXV
b4wBrKU0N57S4U2UBGvWiot6aQQW3yARbLexid2MFpu5DtUPFIkHI1Gul+3fwxcpGzG18XEt6/Dt
HHYKLJ3ErVgPRXfPkOzw6cMDHZU+MMchgbv2zly+nIngym/i11i37Mjb+fQQ27FiIGeuDvB0P/km
P+7yfx/fGa4P6VQ/o/UKiXmUVE4pxZE0DsAV1Z5KG89UYePUgnf8f3NCm2tIdqJau3pWNmW3QwaR
R9CV2Da0jiLqkA/4rvcvpHyDn2H+8YkK2D0Ma/KTQ0LowkwJHVXEm6X6+wdppsj9y6KsC8zBIeZx
XnFZMMSBZhifVV1LIJJhmEVpiMO7b8wSt2eIpeRCN+k91ibWQuURYFZoHTuRTYfKIwTKAnzkLqFU
plUMtPXXLbvKAJ1fRU0JrPD78bYjnBUonQzEx3Gj1DFSNQa9AoPRcunEOioCLwCycKGzgpXvZnox
aP7RsSQxleKRbiZ0HIJxRGpswPF46ko5TxH9pJvcnZGtOsUUvBWlNJVCP5M+jO9P37XXGBY+BsJV
s6i2CxbbWL+PN1YjuG/ajav43DDPXTL2zsh7N+Fyx713HTfi+F7Binooa/Ijfx/uUH/w/qhifrdI
Ptg1wJBh0K8368F5AP7fySVylxoyTdmmPYOt32h1Ys9Vx5VILCOTPs29+oz+GOBXpvOLLX2SXLzU
lb8RHYiAC+Q3XL2hzAwZ+rDZvPfiheHOgVGzVsCgqR/Bqdc6A9+yQvY5R8Wbc6neTbOzQHGV2Nj3
EPbQospIkPlBnABXu8q03rSPf0h97mM7Mgr++cJejv9Lk/LyhrZS2CwB8STSX1cbK9ha2NBV7YAF
9par87oL2UxswFO7Rm8Oyh2iQruvKO7DzGE4CPAGIMBKvzmQqsGhoMpYv7oW1lJLZ9QtHsijURIe
ArIk7dTx3jIpOV50dk1MKrsHT4UUXMlXMuppcBb7OhTpT33XUGDJGyNFTp9gc2wKn1E/Olop6eDs
7EUDiOEJEe93SMt7mFqqp6kr3jISXkeJGA8n+irW2o1EmYa3WVKovk7AboINri9uyGdQpFHxZ2rM
9w+pbvDLyLg4FZrCfCfDm6H2PNhDBzot5Hr3owA/V0N0B00n/liGWf9pQLVX5llAMUyVl27Z1X1x
pFCa24VNclTr5UH9tLr8eHrawQwaMoldhCyopxePiO+EHcSnmZcrqK5A45aDtEboddkS+tBJLjkm
kXA/3+8LObz/XvYHtXMfXBL747YH30b2Lnup5mRMqkiP/XDmc0OvKLQ7BklLzOCTw3dasoGbtrUP
5VMSsK1wihYeiU2up+OHWXw9QUWxTQ5UgPxH80Q7wVKayI1hQJEvn6ZcxvFhZPnoyzJKyfIIi3gX
WXaArEpQp4s0kobHTyiSVNJy3ZAgxWEJDhP6kVx7Z2j5+GZBjC0Xs/MsINz6+j1SlCgw4NTjTLwd
0SOdVNDc7k7EbHC3Peax6S9nZ7QgiMmTbzwiF8UcmupylwDCjMoGaxB4ytmLOzJhAS5iZXum9CTz
w3DiHLo2xuvZpdTtqIryeJ9VCPkfkD1B7u6xkyY2AVNL0d3CQlx8YxLQZwxBrSjccEI54xu4oh/x
OuJeW9CVZaxgY+/01FF3jaWXrnVIyuOkkZDKLU1Hz3hsZQ00uCfm5TYQlns7gn5RIBsYWIJHQmJC
T/AabzQNFzy+O7Q1ENYJ6yadBAquHDfuOr5VznlRYiCyR7fODgDCtm/l6DLfFW0OEakCf+MYzL9F
HHuSMDid5qQn+V1iKpd4U5v/ZjZQrGwO6X0KqeNJHRDbEJsYZzdGzZ/Urn34Wfs322A4l3KAgl3I
JoQ61M5V3NgQKr4l78+LeejVN4V8tIMCGi28BRTzJuD81RNI81tivNk0iLG7znaDVc+uf+PHo9/D
2bxSAPQCmRWZU9ii96vvfLT5vQtJ5lPJCMTjs9rhzqi3Rvu0taVb87g1s18vzR89NyGtKx9P27gs
LFToieLfGPC7/mfcKgHo9Dj2CjSFFnwkSUmFQjW0cvum2PQP/ap12Y2yK30H1+qpYHKPpGB2ho87
LPnq+DJJ9o5eCcnzKUKqiKUJau16uITTW/+Ni7HSZk4tF8ugSCRl403w/nvhjI4njbeIGVRqlQz4
JP8roisKXxntozUd57JLEXSV9W7PZ7DtgsxweNRQ7mbxx+ZquN7RsI9H5tCvvgSbrq6rtP5NFaAQ
1CzimIM4cJl6O1HYQgYxOYMPOqdJGZ6Z5GdgzVLN4g4dJKSxtQgqhKd65Hf2PnHNC6v2ew+se+C8
tBT3hOZ5J2HzUL4uI2WqnbOLZXd4H0p5uthWmbPfYDQ/VrNmBzef2EyYDabjKQCXY6MKcKmW7Cqr
0SkzQ/FwefTkfgmSVctCUGIn4znKCPC3LHQWTWMx7JDWt9ZOgRkjTin0ksaG1W5ks/joDHQxwOSR
m69EYpnxgqVN4vcrZ3M+pB6Q5GYp8CAU+wLAJXYbkG6UMhlov/53F+KipqigvEi1xHmYScSrCcHF
O4C9COq2WQDexC8NlJJRK2Cwpg4NyF1Twep4CGNi1AzGp4xukUO2tEG2+wIYQOAHP2MvC5g7ynsV
nRQWo98tCC9KrYDPH2KFtqcQi7VeSLTp6drpzgrvj244z1J5tGxmA1dwPEkKT6N97GT58md9uPpJ
DSBH2BZgcwUDMTHkXcbknUcaPvfLKS7PiIWDBDa0LhSmsrSUnnp0BkY0d0oA6tITF50iQuZzn73d
VPT52yNeynLxLRyqpH761OhuaXeu2sMkSB6WTTvNaoG8h15g1Y5MR+RyD4iF5urHcObhmHzcuSy+
Vw6MPXRqDs4iQ/NPlB/omtLmPYDasrNFCF56mxtx8jNrxiLR8EfaXt18gc5zqUksvm2DZO7HrXk2
6Wxjg4OzbpMF67aNFpNN7u7R+zInPix8bKUWi4UXgKpcQgvA9fhzZ+HIvx/IRv7fh4JMgntZlIBu
squjJYVdk6s3Bck3d6lO4iFLL9sVEOJxIxSHLOV4T7qV13ylZN+ThKmgPVwTa85rnqBWd1MuDJPR
19apBVT1WGP3WI5t2y9j1yTTcj2m1nJXytaZ7Vf9lhMCu7hZHKECvifeFOsJFInh/4VpkjYluTYx
ewntPZPySuR1u4dr6QUXgkR0hJj5ot9PbI2/tnZMkKRn463PU/8ArbNwGwRFsJlA8ylFQuXq7GGn
95Ma9vT0YdywRgqv4ewJjMkNMG+0jKDkEwNpuCKhfXFy6znVHSjVAxBpBuK/FtmgOd6FhA73yyVx
6Ep1XPiBe8idAM8jlY0TkpOiz/UCQrJRRkzGravQ8ycE78vxfUNwn+blGtdpav1EK3h5Rwho+zlt
BdvNGIM4PQiAWjEWTKxGsaMshgSSO1nCP3rsG6UW4kVHE28oAormIYxaPkkhTX1QY01odcWRWFAR
vJE8INQO3+hmzIkgaPUJ3PRAFvc5IU8x60vjn9DuJ1XRw52QQkAve3f2nP1IIJb7h+6qHgX0pmKz
DxIEzFeGSwfryioLkF41u7RtR8ZjQJkRk29XDytFmnVYkfWHEjvpxmVavEYOB78h11I5/xTTGVoH
knrG//KJt1YMcI29E6IxYIE2le5yMImJB+LzXlauE4sreRjUNJ4bQfX7fqd4WaczEsqToT4E8DqQ
N39tNFyl09OPDaCG5lIcsx8yQh/lvYGRli1PMTznTb5/CaeiWkQu5T9qlpO1dzuniWHoO9oNm9Js
dmxHqEo6NEMOmeA9d2DCLCXwEBwqST6uhLjrXMU6Yp6h4Rco+iYAHKALh+/Mca1GZRBcXRXfuoUy
IUyQqBNyLvxmgw0nl1mhiWFksHnAemVoH9ZsVQrzYPiM8exFJ//Fmt90dUk388cnF0ovP7X/gi0I
IyDeSBV4GunDOfFF8HpuvCrpZrLObRY1V2B7+6oC+IHETY3VYG2g3sFulxPqNibKrr2NECephpR/
PP9bfnQcj+DqV3mKGAnhOOuv0zMkOflKoXxzdLGTLud1z/4kemvdHKSzZweoQAyPcwIXi3azpUIe
12chFoIALUpt4yYCznPt7FLrr45b4CizFmWyn16MQJNdXwv4hySIwyuBDh5hUzzXoQWoreenUk5D
qr6EDD0hSQ5OQrH7Y048AdusiSI1NPdQbpDz2whEOwsj6kvc7skFsGYcqd2+wZKwjUsP2AvRizlf
aoKEl1OIUMIVoYMEqJuT4vCojwOL6vF4jOjtho0ujiNtycxeHcjPuL5NC+uBY++yivoKfYWaqij6
B7854VpKL+RfiuTcjGi7XW5BDqDo+SEuyADWkGR1SwgcJyDxm9YWfFO+/biPoj5D1mnX/7KTYcTt
ia6YtA/pmPLNNsQ8u/Dj67h0GBZgb2EKCWfRiOGpe6l4LRTLI5YXuH5/DQ1Vbv6w6cRdeckZpc7H
W/4Ri3ezON9DLWUrEbsaXUs31dNrTgwHv/oR59pHSIXhfLXd+VeRE2EvKJIDrbxEVp99Jh9y277a
S1Z4MzrZUXditul1lOPImBhEo1jUn19avX28sxnmYOYMdY+RCOxZEasRYXQLSaVKmbsaB23wmnGG
iIE2sx1PR9tFwAqCyAhOev916SDEIgxog9tFuC7UGnhd+rD4ooA2V/pMe9B29R+rwYE+Bt+OKBDe
oDaSlMfhj3qgXYqQxOGunqgS9eKJZpD91vfbPti9HPj71FSFdH+Unz8cy7rRDPxFcK2jKjOptPxA
FMaQgEKDRiJwDorFY5cjbPxLJDKnndyuKb+ImUrO06FV+jyf6TsmkYyO/IIyOkaYqtPW9vqBGsq6
X0HKjIKZESmzEM8bbuhJSuekFDON3nMzCeE2G5i5ydgl9wpRrElJNpLa7U8xNMI2mcPEpILShq37
wYRVTpNv4GSHX4apuXhlQ5/c5NdfdUef4tSkpuclq57UPNGoXCCqyRavv9o6+Jt+VLZeHCgXdkEF
kAl4qgJcv7ExdUMdAv7RCQO1i7HFBW3LbgDDMwRFvUSj/dsgYKNBmtCb0cZhFPaDdDyRcoeLaSUq
Uwp3V51wNzv3Xdbz2jYDm2NyMk2KqXnvrgPT1qVAximuXf9D6qpwCshfVmRd2vCOGrBeVTQwrlhH
VVxHHVycTpICiIp3r0EL0h24kGkw6fr/lOtFT7rKUw3Ko8vAwjXW8SJJgk2yDSpCgtsGHB3+fbaS
zVMvf1OMIoRlzGb1UNJh035yP/d2CxPrYNP/76nmw5sGFQ1kJpQ86d9Bp1YJ9yKT/H8AhBOVkMHQ
DKOJVDF9ynpddLSPGwue+s0CmqtcqiQZSPYFap1y3YTSLg/N+Z4Hs+ogmZCIfsVThUWh2zb75+cU
l/f7cH9m9SuZH6HlfK5c0ZjL1DKcbMz51/hqus2uERQ4jozY1mKQaqlMqoFtFxUzNiDA74nF1Fef
wcHLlObOoaiGsU2/R5ev94TSoT1i8mtoncwKpJvXYZP1Fv9f43lQd4Jh39dNqYe9hkQoQqTMsYH3
VUPtyluSjnOxqi+MDFOXpAPyGMPhk6TB5Kk1vquZD7rQQji6LNc4w1q6Wt0TiuUaZTciqrnMs442
0Dtw6y/i1H1R568TSiXfhShlX9r/6i2O/YJKO8tuYbRUOgrARXNySiRd0e1hZX4i26WQH8tWp2g7
FfONthfJ+1XmQCJGoFug6W67gFHpSFbtltq0BEYd1Fep+1EYaobAhymIvOKVvbLSEqppevKAZpKD
bpEfLLQ+eBGV+ZRjvq/jN9ElIfZ+5dP+SomMM8Dt0An5Oc9zIkiV9TzK8/2rhpVNLPw3djFr9hU8
JZANa0HEwjwYbbwNAWmp6I7fOx2eN9TxxjwuZ0rUDK9/Pb7ADnlquwJUAAM5Uge5NJz6B6RgOhNk
r/FJuhePU5e1SRwts0Mb3yc88lhEzBtizuuuhF6Q/KPBU0HPV95JAIsp7sudXoCPrY6/BB93CDeq
pOxQW7adMm0kc5E45DAAOdITbWfso+cstUQXoSVqukv4OWktxD83z61M2s09rm08roKpUVBi16cj
TJSVj8n/QEDg//G1mWy6MnPCDk0XHWzAjZe000AJZxp3xlHhhaE81t1/dVm0Wbb6KIUtPngt9BbL
2PcIE3nJoJ3+rxHUvYXVDYIdo6qWu4X6SysnDoRFw+KEE5MpyNftGHrpUeNlPv8eGhYJGukXIW0L
781PCrCx0T5ZYuaG8G847K/3pTplmjA6IiFJHYROiJIu9WOok4WydSOItkkJgmxVf9OMWaTXNtfa
/1MXedSElc3B8ErMEVOSQ3D1i20yMkejB18yVYDY5Zro5ph22mNDh5CFZUwVquW8Mwm6d6aZ+yKK
NvV0TazNq/yob6lEHj1xCRbAlnFiRyH8aWK0qFzVfDv1bJPA0FI1P/X7Uc3zeI1y38sBxuvivvyy
DUopT++G7814yZL4p9YX8EV/FB/E1PX2TL2J5eYmD5l7UM426+ebL9H7GcHNxe5ADjI5BEG3Wtnl
3n9+ZqMrlvnjCWGcbcv+t6lspFycx/SARlf5BdBzSR2niejRGI26BbPwVGipQihKZ7s8SiuzvLWG
hw8CW6+3rURxK5DNzo25fUyQ+GNLu1521Qy7AP3WjglF31ndngLeIHdIQby5VtwOaAlTLNFla5tu
ZPn7C3WX6mdR+GeoJwYTwjuTWN7IsakZISE9ZWAFODDsTVKwjYFw2ALmaCp0IJr/tHtdaQu4tmU3
U68ZbEyOQac0aD42GuwGanbtyySIt5Bp/g/RinwnRVNjkKZaWqIa7z5JL95+q7x/LgAjGm4mHJZe
tXliyzcw+fPpl+jy2Q+zghwJ7hQMr2Zzttfal+eqTyYTN09HgIogtb9HPsUWTudVtIX66ju1jSH/
rdYqlz84GBtJZw15bT5UQ/94CI8gg898V+W4w523W1YYtKsn92EIwdvMdn/rRgrmhsG+qGJTPoMM
9MaBR64MlT/4KaTQxaESotRA7Tq6hbZuEPFwscdZzbNp3bHdQF1qZ+M5/nzjh43RCR+pW/vEraxi
O2cMSenQFTS+5kqos8qMExejn8gKjbAng4IjDtwPPUKvusJRGYr2eHuPi7VKIBK/IaI8Z8hcysfR
iMeF7Y1lIslQ15eVGJ3t9NgvI4XnRcRyBrG/4/ctvwIaS3HEdth2gw3VGulxmFoDOgUd8up+gHR4
CUqg3tU9CUwgRXU3Ko7sYnmW9dewU6vmV66dozw6qWbS6qmyvtnP/0ClOUlbdXnyaAGF7dapxFDD
rdR/lVCFzCG8a1pyk4iu5hn3tf8AllJyMCviJkCCtNpuCylEoM4w4HYZK+sUXmdnoQkhAGjailnG
L6YmFr809umbdWvnfx35XmNLfYHVkJMTPrVjTCuoJtc25fITTXpYHqsGcCmVZgAQTehQs1BeIos4
CzN+lvqbRsvf34K4g0OZ4JfyoeIszvnTJgWVuj8zAWEutsUaDSfRX0GXPwbFig/+fR6hSsJhTGI1
PIBnl0Xgk0ZS0g0gy2SwvmSm4qKv4G8oq+ILvyEN2CH0eja6TO9UqvWXmPXMUwvKobrIeGzIYC2C
WblMOcWabl6fmcJkv9kmapxLgA5ogy7Vhqb254FjYFXYz9R2XlEUrjOzabj+0Kd/WUyCpLGEbDMg
yC054sCsZXrmomKPgpUxH04sM8cej2VyEhzVOX1SC3g/GAQOoYH+vsejzKiD5EXHR0u614a/DXQ5
tb1pIHes2yM4fFJI7/lYQ8MJiXAZqKIMCNkk/iK+paza3ZhVnn95OOh536D8xYV/ySSXeB65bnR7
ORA8jlN4FGN9wmdtgyOKqEcI4iTvDJhKrp9JRKJwinNFT6VNx/ZeTmAV7Lad9dA8dTxGQ0wkBbfQ
Ne/OAdQbZRiXyMF1wAODofsiYy+EknIPe18pvDKxLlAvWBHDtlSQOiK6PBOcjMrNyvgnxbJiD/lo
ChmPa+TuPEqLZWJ60CbYFl2H7i6dGFpw0ZRnNdFcff3CRyNs6m6HfhL0RHDcagZWxIAdTKgEOhlg
A9Qh5L42/ABPe920o/MoYskT7LJ/t6kakEDpsGf5J5t34hWfj0IIsolPz03OXGcNETW2FdL0zA0m
7VfmlvQHjfjy38RI98fRYiEG9T2/BuUfpjY3h/upIclyDrCDX/GdPUdvlaYmybWyXkX8bqckVhqA
MrxGF4jwwpRtFeSv3N0vii6IxtXeGmanfwrTdSVhDe5nSm9XsVYU17RIvNn0D7hngxPzwx2+SnnI
eWy0L3M+L5qeu52TS+SYq7vatvN6y6Idfc/uZz2VzqlEXd1QJTNvSrKmhwMOVwmvMtBnIKy4juP6
19oT97ED6QQ09rekdb69FGLWlDQ5WBJTu/nUR2L97LmiNZrutVyfNOTpyTMRneRwDSHqeCSCzgjR
gQWthyzXWMqwzlu6y3DFFJ4zjATjD4PfayzdGBHjwW+EofEPS7a6LxJxPN3Zp1jv5AHBGmuV6pfV
zKs68iX7Qa/a74spGA46lF369cDTzQn4PHNoglIeV8qO7dga2RqH5oyFETSeN30e4iUY/cTO27hQ
PhT+6irZIpBXpbRQo8oj3MZjgDhtaRNf3a8IJdD2THuaZanrafjMXo5Ab3dhhf3Jc89qotsvZi+m
RU4LuGH/ioYqsqW9m8Mx0zvHTdMinL8wjCXZ27Q6/ZfeqNIXqiXNCXz1qFDVMMoadGxdSbmkV7d7
wWGJNiOx/mA+k65A/L3yG0HJDBjoQvV8A3YgFtxyMKODCXbChZQHoUgE5qAFovVp7iczZOPf9oWv
609n8sdMw6jRn9xydKFyL+sH4VbsgjC1KcGrYSuGSNOPU37A8fLN3segOb+noCg4ZFbBJhqrCcT2
oQ9Gr8dhu349VapEUh1jJHyt4ZKoh5v/WviwvGWbEXS4wjJABBlVEypdy2JX0Op1eNGobhCqtFma
E3EFFz9Dxx8yIkVqjH8PzI2FBHD3E7kmudL7dm7CUniALZEHmRDyZvapsSsU4DdTxeYGMUfB6PbT
usT9O9LfpbqTQjCIBycoPOc4ysVWDl4b91LJraNeuFrILmpe7t+4NfHLncV9Zl4m7X7ShqGBQY4t
bB6NyIF3RpQp8STjcM0uyh+9oYmO1ocjHtcHjq34XpfAbe1D4QAU9T/NBmKK41K69VNvrJ2Qkmhi
mwv3KfKLbFTUfZB/mrjR6/32mQ4fVd+djOYJYnEJgJH2zZQJDE+Fgm2Gvq2cRznSPgJ3TYT4e8Au
oKoatBdUmIEdHJDoAqxVR5fV0z3j76gMuuAIoCQcRT/kOQ7ZfvxJ4awCNitVSa/aCZOECCUMyQA3
cIh0tb8ZW2UgnoIMEWrr8kb2dHr+2C5n1ZxGhs775lIJWYop7/3ouOmhy9A37LFAUIuDGayeEtDr
GfDgRKLY2l6xHV0QNRkszF6rsLYLudajQ65r8yGs0/8vD6PpfsEliy7IhlwPlSYnx/yzHaAdBY2F
175ev2J5QNf7WFiBmx2HqfXo9jxLku95jmeg+XE957bNa3rjEr+OWzghK+PKAKIqIBwFdarPd0Dc
FY4fAowlMpD6Ds95H17a/ctEI+K8AFmV9nH/HFGM5X9wdXwMO1G0+Z2k0ytuAkW88qE1H9KtF6vm
TNN6wImynzeGYfjjyGMS/ZKpCsE8FNwzO+0ajx/9rXD58fb1tBlLpsHBWwDSosaSSuUWK3JDqH4U
Hyf50zbs33+GmWDu48oufq0IY504fHp05yNCwfcdRiSgo3Z1iK/Ohk/4gQT8Tp9XOUhzo8twIzys
yMybg99JdAqTef7GcDKUyDggeZtPu9RsYkuL1WckPgMNUCv3O8RHEIspOSmD6NoorbeqLUYhc6b2
BGVOka2IWd3o2aPnkV97bDtbuSK1DH/amNJ5JBkqhot1Nc2ihRPefKRF8KwAglU5zws/MpbzFOSk
mEOxZ+Lg3CP6TqrBbk5xFpJi42LVOTLvtgbl1hRNYMV52AHrvME8x5lfo+GB5Stfvb8QxdS/KikM
WOG6apYAaEchkI1B6C2DvxwALlkgJEGFkx8qMRgRcHrExFHbT1tF+dc4oedv3U53zdOzDjH0iiD5
iu10vxCsmASqQ7m+Qqj6pYWSCrP3sUhBhiPp+atratDI7uOPe+gVTtIr3bgSlH8pBBjkrEgYl7X6
u7tA9Gp9BTdMeJKQJi1n+vDAzzJ9Vud2bR3IbReGI9ONqYsw1vcc86JSkD5J/8L871HiJMOo7+6f
xky6D3ScDaXx/UFw/Cj5JkFiyGID1pzHQb17S3Wa5M0jObyiX/8UuuMaW7JAQ0zlLgeLVw+nFQFW
+otoDUochkP5rYK4nNuKIG3/RMdUmi4rr90KH1i4LJCv4SdnK7ZCJb3W0frsKcWSNf9513OPRppU
mRktHBd7VjOVMVw1a4oJovD63nAfrLjFmgOaIDggONIPVZ0/kwzFs6uUy/ypnKqKdZ+9zuj0Wmpw
+xsjRV7zlNyrzbt48JUhu8ZQh4478iv++oZ0augpzhvIbTm8RByQz18vb9PZgkEsMiIuB/d1XK3k
30jTew0PXODdcifGT18weDnsUZg4Ip1n+177R+hFgjw7vGFLxOza6xkD8tmh2R1Qn6jWehPnB00d
H+DcFEiUzoSUpl95E337OFBgrWo5aFbUbrZFQa2dqWPVRnapB8+N4hCbNJi0Yxz7UGeiPL7ybfMj
JCV2llJ+uPuw0s0mCtly+rGPtB352QY3mSYqi0kyMDC/sEQfhtqWLoJqiyf2ejyMPrfvHdbmosmg
7LxJggg7KJfSTxxF6x917yyCn4BvkXRSogAzbFgQIj5xb63daglHfOo5KHmJ90jB2KOSvHVCihAO
u2rMPvXGSjxdB9WkZ61yzWJ5IJvIZ7DTkxlwuoQgqFoswM6qX0WaAESsksxdMbWgiG0ic4Um2Ibw
kieYzearzd1rYCtWcLPwIBaGQiUl4VNnb74Vk7esXCZW9uJGxUpHLnMCAY0hN/KwrIwu+xVz8uTm
kQKFZ6wETfGsvpHROzV5W2kO4VzApVrQlhfh+yIQN81w709LNDMSrsQBqJzlaKj2HrhLQCka18IC
h/H9i1uMBrmegUvTq/Nsb9sSXXTzfkP8QfZUXUzFngB+DPE3QDZkxQKIjrk1BWYxl9ydLFOkhXaT
+pjNJerTGfDcZcioycW6u/S0f69Cmohh1UCLeaD17eq/PQHTzJ/qNgyuvRkMK7iO8BtGrHqhZjHB
A94Wi7J0/QoyTCjRlCbSBF9Dv0wO51MvjOEo8zBDWgd7t5W6a+jaK7wFg4xe8cgb1hRvMwMfatPC
Orq5ku0WqySfNi4bPEv6gc249Dr6+LixI4GzojJL/a6C+tpLfQER1AStZdbnhnwP+0E9S/W0Rgzf
GYcQLBUo9f37UmaaOTwg2vdvR5sOCG1p9OSMkg0xbNU+beqUFz77nq9izYHm8F/qdQUs/P7cn5d4
wHOw/DfLRiEBrO61G9Y9petdl+yDsiKulA98HCewhAzf/ePLEF/OTMHc5dIYOQR7aYJKJ+T4psIH
znenJ3Q2HNjtNmXdtc0sGbzVZE1Q8IvEaL8SIKdyKexu1DwBBtyR/xVUluJEErPORl23q5j76RYX
IPjXuFsj/cF36x3RTvT5xKPPZss6LNgAUjF3nUC4JWI6d/17HHhbbM0j6Qqi553geqVWVSU+35iv
XiM+1NLTrsR4o3uDS7R2yAWMq5b+KKE9HAARIQgxOZmP5ts7idoZt4F3HzO0zY7g/l3j9k8VcQ7l
XlWblLEobutIxUB8TFh3qg2rp4AiqVFiHW6JcMnsehwbKhQO5MLJ5xPOErY7ykjxkcwAaYEpgz/+
7SU7UKNOTl5H2PtMkNkli8oTn7O9cvIMzXxsLXSEQLNughGUrRDOqpoyY67SO0Z59+7DwBcTn1+p
fZmJBq2sDgHbGpI4esqiXYtKapxSj01gti/iNt15VHq7q08uzgIeyHlrH/V7VVrusGKc8sBe2pvi
WiqzqFu1ttiWxSKwKXUTL1bFnFLEpUYhNAANdnDv95NJKpphBa14etwNmVkVvDPJi+hPjQuVGcbA
vf/GGkc+L6DL3MKOSOQKXtSo6b5cT82kvofkrp3BMrhOGpzJhc3Ryz8dgOsBcM1gRrubk0H7Wrcn
iO6v5ZWFT3tO8blyCjZNo8DV5RLYUni9dKRHQL4fQC0BqlXvTL7Uq27NY6grnrSImBWsEdAFxhe0
r0VJuOjByX7L/Zcrhzk+Mnlp2Aq+iEPASQpKpQDcpZzqQHwINlBHgsQMTMK/u/juoq6xzd9XVAI5
oZmAbACM2kxgXM1vJQ+6xrtUInr0qJgpWuLQtEiSnxK1KQ/y3Z0cwELlWyNEXrMeEdFuuk4xqofp
8p/4mnRIVDTPOKEh0GeVgGzUwfGgsNwUVo/8KiPpMdTA4MWo4e7JpuppGi/glh7Xw2rOBr9Bndw7
2wDg1zYaOqljoyy/p1wvarTg1lFvkzoJhClOL4dFumSj5iZ4PvVU4gJX2zgyUDYit/hOtXGUVGEp
TupYlg3SBSyb2UbTHJtm3xN64h1ez3GtVL3JxeWyvs2dvKGXSc4Cm6o88viMfEb63RdM8eojcXw6
7N5rwRkkKDrjXD9G2NQV1Q0D6zHvOAohhMerRpZQ7qZ+xRjMjBQef8I6KzuaWIX+oZyq+1bmZ91T
Nywl9gDwSsH/Sb05018DAfwSe2+O2LqAiTP3GkOA9Sj3T5pu/nTg5B1Vz2MoT4yme+m2nJ612d3h
ctKt52XgtaUn4PJFOgL9Ew99EJmoKKQoGu7yOlSTB+Dc+VdAys42tQNDEI4Rld8Rzx6/f18yB8qJ
yPeROWihAOajs+1cL4stKGEI/pkL8I8qBFH09ZL3nWYxpR69MCb9DUUcsZSq4hOnuPlt2gSdgVm5
dwvAgXYz6S8dgEQSegDdpXEWpqbj0PKvFeXWLTVwwrDAPVdX6IG6kl4j+M1/tvGCTykyaoHf9jPl
OjtWvc46kyskL+WHQpH9ajrBhY8eQkf7x3GmxrOg8XIQHv2ojLoVEgJBMrndbajk/xkpbwd0EiJb
AxATc1YfzuqTfKN59aBXaNGY5dyR2TzPa4kjZMtaJU+NV7lIaDSzFWAeI+rw5XjKpBrRSKoXEJ50
S0wQvjFipeRyWf1ulf1/20oCv3w/MDZAxSYHcaijWOdboQRXwfUXbHB1w7NUb+h+DzP8pUNxhKV+
LdApB5zlt8FNK0FeFlQRjjwif6Yc8yVUh8DtYh53Hl75SwOVmu10Udl1b1tXtjcszohyHhDWuN3O
1RILUuvDKvSkvKaGboXcv7UgShNrXCkQj9t7/57fU21GuWAxrJEX2sRcisAsAKyGKcD09yeTTXQr
u0C+BOvPvFVqAOQwmrtFQqZ0ioOCadvZ8sI0PtRUlFBPZJWy7bHR1Lb0pv71mosSjjjX5+/iREGW
FaFAuEN9q/wbGpL4ZAU+0PcniJ/WHgmUGz+q8xaTizZBKkFVs2xkTnw82DXZ1qDO5oqwD06l4HV7
tRDxQwc+a7TWlcXcDK260LDYaakzl7gb+ykjmJsliA+NRjCTzLtfJFBgXRRVEtMARw9lNBuKGzER
NoYMrP/wMTJZYPji7m0jt5ILJ7J/jGF2AaKjJAMVa5bMaUS7jZw/GN/mZUn4bJL9AS8UtTomG5ol
TkUhKwBcCIt0XpyvaHZ8ifwe0l94LI4pwtlXg8qHUOkVzqCIrykDh5d3YliZ9LPuVFE7mugmMJnU
dm6EU1tbu3SPnQdYQHkfHTwHg4tqpm98E5Z5e6H3rLUGTYuqVg311fZ2o6OR2clDXK/+4VIo9pOm
Eix49HjhtLy85UKwgRRZ0PO0GTK6cZnLv5KuimlxGcZhzVzi6IsWHeZGFbsTLpyLviPMdtOtDekt
pCXvU8AD2ZqBIlAbAAI6+ViM7M5Q1jTa+h+mD+bHCTJIkqHpbAEDE95SbGIV6koskXbz5CpZho83
T8Xuc7z0hStwAxX2x0XfrWoTkwQjZeSO86LuAUEzIBdE4NQccmIB9qS7Jt8NtajV6n8dp413KSNR
J1pY841RPXPe6aW2xdp7VtqXyYqqUqQYCaCxf6QbTfae0lOwaCCKb15COrVjDa1kzSkLCNgnnh/Q
0KdWWEjDPJBmdc+c8Z5esrH4+S2iwO19xst8jZS3Sp5mSNWCNtICZReoRafrTSmY38CxYxL5B+n+
vW4ocGR7t3UWqvWE6YV2LJEi1KQlimhtt+zNKbxwsGa458QXmXNNq5D6hLh7UMAFFF6AUtF7eTcG
N2nWxHr8G+SGC2NtXA6XOfcY3+sf9gbBoiIiB9hl6IWojANWG4CTHrCSXKBVwsRuPLfLS5nFEjtS
ID+cH7EGY5gbP29AcBohNVG3mnu0/GOhu2zBZ2llTvW1GiXrztdl8vQrPxO/HYC8xq50Z6Nftvz9
Ls9EDuU8tp6jEUyZ5b/Ha2WMGLKW3sw+B24fzz8UaE4bwJm5sXuNj5a6x+beYXUjM/ULDEhg5T8s
4swF8Ms+ObrFRhlY+HatQWDV75vmwSbZ12QJKFhw3uDmKgqAxCB6X9imYp0o5wxnIJ1BW87ylcIK
1+sp+io5BRW43rvhfXcsh/OFus46L1NjAzc1ss2HOs0RLmZGxT7s5NtVYwN6D0sofD31HWQLaolX
+HCVq7xl5PywNpf8gl9F+fuaz3QX1pzHj+7ygQIHYBoSZRusqk9gLtaorcZV0fD19lRioC0fXT8F
Kptq2S5q5F5RHMUnEuy2lKIJECA2Ra2l/PmDBu8Jxfv2+mX4WVhC9L1CCcazP8qZeU6BBbVSuVd5
GLvVkrTTYqwGCVs3cYqOMv54QeNUQWgF1xvmTWaeS2e9wiYg6nLEZSlU2sAy8EMiUmFIZMYmjWz7
IG2H7FpyvtUG+jzx06H85a3WOa8JlYu+eIlDFkNzpKByagkvcAFm2Srbva1WA4Hcd+5Af32aaZZ9
33X7ooxcmsAdPZd4SwFpCi6tjbMI47HUuf/nXW9xb8jrBlyuTq2U/5A++KkT0RSsHEdmEXO3wXe2
RK7S0X/AnqQq0GWUouqR/6FSyNijMCgVosLa7rEKlwqADEEnukRvs4Z2LIqfkwSY4JFhF2lSyahc
lCgbk7RQ9hW2igzowClhshJdZHomag5E9cLyXV10p1Is16Odz8LCqQ4mrHmCmPB4unjZWV4x/9mF
BtXBMWcn1yaj6TxnfUusrDzAt+Uwl8Hkl15K2Xxouot4cRmXddFOE19nYf9X60XxXdK3gl0MHzgE
+SpTBKCLEHm0ooH6ttgD0nHAoOsGfxX9ROFcisEWaMLjMq33nKhc7d4BtH5Yubj4cJgMN2PU9Tzq
lSkvWONYvfG2hkUU8Z+nzMm2hPvIiKyDGFgUHePBkaaTzkl6AWCLCW7kcXretkszsUuoYb2qK17g
Tytb524YzE8J/6cy62MmRVKS0bwlQCbOk0jMMVTBFcuRwAZFm+zRkq4oT/Pjw2eTUFM67ZFFo6nH
vxm8SV3PvEidGJz2b54te3KkS9CIj5YNRnY3kwjxCp1Rm1v85TJJZmDhxKkKyQqFmvMB2FxWI6gY
pdnOGrqSPFm5WdWidk7QDUrcQrfBmFLOUdvNKnlesfoyJIaB1kiGf/YmHTUWW5vYCeiJphg02Eiv
Lm54EZTmcmsHAy8NeDSMdgvvQ5buEB2fWynr50EgfCdvExyhKy4Duf3CEL0qZk0SOq77KvEEd5SU
PbUQRtuoF0gmifrMiKpGsrlI7j+4yin1qPZhRlannvpfzamHYYt5mUU1QYkzZvA6UCkTCd0vcnvo
q9hyEA7cWoFa7y/xkiyuNZUx372L9cHoCi8Xc+5gixkytw+aHFNVdYvxAHG3sRBwFqadvFO3Q7Yh
3iaYLmTADxR6WG84iDbiWybu65TCAWwYcwFl3KiIpM2H2qYZpIYDrKVBBU6+OFGHEdntqiRHlOBH
57Ca5a26BzQMMcfEYYGKrBp7HF8gkk5SBs3sx1r0yPW8uzh915sTwb7b6MOc3IdxtnzfgF2lbkUT
kD40MGDNpv27fjLQZrtX/R5+Ac6JkiRIVaJiFdDQxYzsd4WE7lztyjr0CTy6nJ/cOQmQHTOLmSS7
yNjni9dAn38Qc/AL9VbFr5x0hzoETe1oJrRqj6f5KM1h3IqhBvi9QNk25SN/Af1OGEeaseEiS3P2
ObLdnAf4d/4xlle/6YeTC78XDlec7JvTcOr7EjRiamh3Nm8YS9xL9EINyeD+j7Sf+55XtAsftYCS
0Eujmx0QCy6qZj5oaDZPwqqA6nxj6P+TSUr2+GGv0HHDTPlomJMffF5aPH6fg9ba6jDXInvgcLA+
gF5EmQKDcgCrputqMacvNtBuv+qe5JbgAXJcHPQ089+mjqRjVN4PuhBSf2ELWw/z5GTdkGqO+Ave
sgDMrx+se1K6i2Vt3dO/Vm5hZx06fUXDO91qOYIXIJn6fmjQTSmNhvZ9R85HntiUJFD3VeXPPACU
rsZwged4agFYdm0lqIRgagFSpx+NXm4vYOOF9PGxJqsfVCKGfGGM81oLqflCLQCnGh/fSraveesl
nrgOn73bKNhFv+tagKC/d8iux0+SKO1KcQq4Jp1tPDPwGioWmvr68fsURFzMzirPGIP0oUmpcLHX
ovHrcSxgME0L8WqCTUpNJqKaQWh5qZWrJ5UDqIegYSpFnSLRfllvHbGdFWCtyW9tuhKaJOzS42+F
6/rehxE4tqEoi2gT5hbe+8ommkMXYWEEWEDQ2rCHCbBUMLP8yJoXuzQVg5P7nIeMm3f5xr9H2yNX
rnLQ3PgrlC1o9aFceMtfEzxyL2VXaaRGlRY5Z2Vrj2YfRX06flQejX9Bjine/4+zT+r2n+WhW0+E
0XXPB6DSxVomRx+6r+96d/89MxDw3bxlXJtUBHrhqf7SvL0P+SeJOMpq+AR3PBz3dR70IePRz5uT
T/avzw3m2yAuA0OSe08dC9n6GJ8arjpPTmNmEt3YCBNSqHGr5+HZHDS+XTqwmsSFaDnT+DBlgbCe
WtmGPxFWyu/Io5+FHL/duNcgqDoJ0KFCGPs0ENs4TNJmPRkiPTZblMmcdPWyvMhCqCdP6MPK+jL4
7EOLPM/yYLJ+WRpqGt7XqIEdff5tO5gj2n8yIyJmPHlHunOGiHSBcSdDtgxpkHT60SMnEfS6qwn9
D5uxMlQh4E2Z6bY=
`protect end_protected
