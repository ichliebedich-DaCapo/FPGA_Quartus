-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
U+vj4dBAHlOut/dBAQco7aP72tnKwGJgShmKlhKMaCPh80NqKMal2jtq7GkYb1kV0M1J9HvszIYL
lDMGVGUBCTnNruFUi4llZIEEpLHmB4O1Z69XLIyGcagCZSI7Mcmi0hlJT1iYv8wKUlonZ3xv54/6
P1pL+xGEG56OZ/VUdvwV/zLcn+pPJtsWDjsGHOY4zizoIBsgxIScKKxHQL4ABRkpgTfjt1oZkwkj
6LRDMqz8JhUWeJD4SQkmW1klHNtSOLUs+NDAaU9giZX7ahITnT3yu5bojIBn8Kw2BRhONhSbL8x/
bJbr7AzzoEDbQgv6cZELCRd6IIsFQLshOWa+Ww==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51056)
`protect data_block
8R2eHtLVwt6EZDShw/8HGW2O43j+USrnKd3elFBDxmSH3PFvZo9xurpT/JiC8wGJZgmNIE6leIDP
ooFZqXEjnN2y84stMvW1wLqgPyhtSYhT8Sbp8X4taCQIpLPtoIRDIrnGKXASbWAjk/8dq9DpOFsE
eqfbvjNZ+SSBjdubUSEW8A1eXBEiMwK+3DlDWzoqpZXGKUg7rKVRI1IKgff31vtdKjjC7w+36EEw
zzWrTpRPXCnwku2p+0GlH3UgW1HPKodnoFhuF0aQ1/td7NLKzlZTtAb6RmwWq2oQOM195xfqEhB/
5+0IV9UzxSIYWf44mmKdIhFzL9rE4jsyqt2C76JZZd//cawQxF3r7Zvg8HFXxqJ6EyITBZbxYdeA
t/PklqYOBNxA8+djG3JXSU1HGI9HnKyBJeg9CaA9STxzZOP9+jZ5RedHAUqGTzFfHLBllBMu0wH8
WlmWHBohc4CZubpB0KkcQ6CPPz/fwkuHEUgW8b7GzQl0K4kgCTd4Sy6BO016c89D3EjXpsm08vah
3tX26OzST64LFujRo+oHh7DLsO7Qz07FGKK6fPpoY0iDwxBOhFV18OTjmF+Y9buwpDUPFFWqmLpu
sY0fQpq4uAhgMp+X07kSTp8N3FwyvDW0tsKZkDSCu1wzuUqFjTrxmxydtqbnxtSIZKT1Kl+zJNMt
0RWP6EX14Vd1FRQqfU1mBELT8t8r1bp/xgSzpCVtmRiaYZgnFzncZV+GdNKCxwfGywlFfCs2q0C5
eWrPTkJ1R0OGZ9tOVwtWMYVF/Fh+zkzf7Zh2Tvnr9kdSV9CwsC7vHIAZTGxYhszr0tunHhw8UwhC
qxaEg29gASvk0GfHe6DytYb9P+hSTyCdsY3erR5ZBEqQmaGuDape8nODMx7q8sijH4dpcKPQTghy
EsWjcHqlUo8X3vvHB5ecOmaxi/4L5voGA4OUL6povO+7AkM/n1rhHZvomJZ6tqGEXM+t6w/c6xsW
2ivZvJYPnpJegYthG8DL9nSCgScPgv+suK7aJ7eCcyV6Brqp6nVklQu8pbPz9SKiCCihYn6SsnTG
apPPgRB8xKJWv0CUOQgdTLK2szWCGpDRnER0bEwHlUZtsSqTje/mNLrjhQDKVoQwlaPBfFSTvxWM
4M0OI02xacVRfM/9NzHZP++F1DdjR59Wdu5H8dhhWIBSlfTEGP7xpY5VvbM2RRJdjd+5RHisB0XB
C/L2I37O8gVSdjUEwC+N+ftt5sBK2wc2ubSFDBZVNNdL9D1KmA1F7w6z+7azqroJd02xeH+c2eQd
E+bKH6VUzH1vmw8M8t4Z5UkE/80elRCRGRqKy/TleisYf0eva5RpG97iF/PiLjiLpQx8Bsze4mbc
VoM8qGCEovWhBP1g/CofkBMYCHVPaLaB5qJiLoCXB6u+A4hdK/iZEwd6b9ujS3PNw28bdNxnNhNx
w1i4sW0rkYJmlc315Ul9ZqzqdP0A8k6dThfXzmWmjn7Pd5ghOokNw0A2WTT9hYJbAYCVTdHGJlT2
DFbwu3VpPEkzhI8+QSSX0ZZPDzhOuCKlPGsdCBoGxDu/UYBMYNvyT2Bs/CD+uL8a3sEwrhMR9clQ
fwEDVSVsCAAUr2MDG3LdfZmX8LOajMxbD0DCMayut4bDYX55NJbD4yrr+cFRKb8Wt152u5XyvSdQ
PPc5Z5bO8jeWSLTHUyZOlVKkXkYlyigj90LJgiA6jJ5PQGAqMzwzD6BtVEvFfI6aOXyJHguilNzi
RnzW4QrYRe0DFyTq1o3p7B5sRkPcpAOqPT89DI9nbdxP9jFRH3jo1YORRgU6fcatOVJipA3BWreD
e3CClrsBPt7NaIzSaf/4OQUYqlvb/kVb1gDwPFNaV8fFqjTBhxqyoOaEBDatrMAdkFm5I8XBvDI5
9Mgvaetypt/MzgXd9PJ+ajFSFZb5CPBPnF6LnfS1f3YaZmQoFSJtirS/ABa4m6EphH8C2Fhgc3a2
sN1nqeMaovJWAyC5ZBP7+mwaOL3yh+41mwyhivuZJfZDkwon3AdEVwLgre3I6bmVBvCaBZo2aw99
zUvGb9UUkTzr8YuLvZZQHxmI0ILq7s83cL3tuTb364NrJfX8hLQssmXmCaKXkRMW0+gAkoRfa1kj
Vs1c+pUCk0p2bX4mvXVF27usNNP/q1PfE0Y8TPsF0SrNe3H8Y6w40ginIc2g2kIQD79TT9NrphiA
U15WAAalXEz4JCpJz1DXFjf2QqHnpzfwUEKZDG4u3RkPH+gpiubmFvuA0EOlpoOq75GMTt7nR/Ud
5UlDTRoQAKveUFeR6/zkybY7QynuqQW56FEijHXrAB39lN+cFc+nmb8HlniqGclVwaWcVwF9MTWJ
r7uNWVjTnRnp6DKzaT7/1FcNvo0EPgT7RC9WRRODwsqyKNfJq0WHebnO+6kYaMDkE/S/q/Y6qwbV
Ly23hLkCautx/Fbq3Um7Kje/qw9zC6GVajPrTRaeA7S0ZcZDk5C4PVUFvz21OaLJB453CiSAIG9V
oK3RuxHbhIEIdLh6QW8QdunFsQUItyOy69KT1RAEbe8D1MDokM7CHeh6zJNQZ93F9zyX8eLa1qiM
VFKYdAX5LWTNYvFcx3GmCJvGjjzZHa07E/skOClWRVpfE4isLq7e2XxOv9miQpGwJxDSQHNUdGYh
He/wz8p5e5qV2YC5n9pCUyHQ+RiXuRCRtVtMDnIj8VA9OHSyeT1CR+I18bPyTzXX7wrJhDrxC5Ar
x//SZRTY/ms6u2yk0ATt5wQPG5u3dE2syyas3xh4xQ7p0a8IPwyD3h6w/7EJy2iVmWBD3bgGx8F5
QZjgqglwWIZIplA7Z7MM1QSNcRGmhp1K7HEl+uxeWx5Y9Ke/69/kQcQq/u/VdD0kau9QV11IP+Be
rGKw8WwsBH0ormLloq4mZi5C6DbRs1pLKI/H67lUQpCK5V/VJq7mu+jZe24ckbHEpcEGL4i9Yypy
QLpCG95GJsi8xppJkzt4JPz9B5eeslHeeaVGLp8X3MgovXczCd8P6iAs+w5wWDIpOd96eDWdB27z
GCIN52Wk23ixo9uWqR/vaaswYwyct4GfCzIGi6kpO4/Jh1KUm3l61J1BF+ejEvFn/FJ42uixkm+F
SuPhVTVgPmZcO3UXGLO6ZBu2GVThv5pvtCGKxa8uXyEF40PAKqRL5tP0jpR/te5/Fcz11gq+YJCR
q9eQoI54zcuwErC3jN+Rv2CmnhUxC8R+IcMvbTpTamy981wCuIO8mGw/UxZxTlY7DWMwIlxLmI7M
Hm/NK3wd56qckV5VFCCs36z8HMBFkUIO9xfpyv/k7T14G02GDSHjZQvVp4OrGrJN3+iVw+ESFDJ6
sBJjjoNYv51YVwZTezWBtE8v/Ptiz3bfODXNC47c6GwMfj5ng1I5zhcofAWoSwS1iUZOZkRbOSCY
X8iIaLvO32QGfjRsVIZKyByceChMbyF4mYQ4W0dEREHPCTQcwxB0Tx2Rh+r6YcOpXzng8lk6Y5tc
qJdeZEhT97KLNOqIeahOXdx0C0X9ZgVd0xTTJ85q9VNLDamtJWm3pD4hFE9/ieTcWCBlnPtsdvY5
jGvFv1wol5YdluhyPESrTsLtwfyEV/hjBEiczwuOHZNVj24dCzsIVw9SreaiRyM2rmA+6GgujDOT
Xc5WxcwR3JXYJtm2J4plq5d1LcDpgoYCu7Gcp5hJc8zYvZpubKdnvPVTlIzVDFos/u+whhbkIq5a
y5XgP8C/M1hL1lidyh29yYp4GG2z4YQythr3gC6kwLZaybVpQLW02jSq5BhBScsHUwZqzJ6VIjc7
xudP1GUcodSXogYTyQ4unavi4JdwLA/IbnGiB9kNOFxaBn/eN9VKy/zrXGjAP1fM+M4xV+SG7sCO
9Om1RyW2SksWNlRq1cUUunwVd8E55JgF8KwozfQPA0XDXgR9Ex4j7+NBQP2GotgMxs4w0Kv9QiPH
FnIgPNKnhT5xJQx5clgRVJuAOP+DnKL0uIyqxEPtnzLqhhj9b+AKjq0k5YSjDhtFsX3VVdNUqYSQ
Ct7yAPx+9avfsGZWXhLiVdRS5FfBFqataIq9Ts2uSVBUq4Xywz0pBKK/zhIJdGbwA4o8NPsS3yWr
tHnH1N9inCXsNL1EG4d+6ZrBy59AQA/QT+jWPAouR6Do6zFfCN+l3XOhWXqwaqCyTFuYF3EPVoFw
1EBt4/hls897Y04mamVt1VrrqIYY8TTh0pGBhlxJu1DJP/KIPAGn4N7Q67rpf7e6vTmCr2nA4qzL
GGQwPz9lKb5U3W6WK9rmuoTBL8g/fXAd1CQXjqInAjJjXJ/bqlyNKENex5So7LcgUTH90dqxhLJa
ArAaiCGFOIFBXEdQz5O/To+YIFkOGGniBh8Pel7ZD8jio9ajp0mSB29jJ0RIlWlxqcpOixCRPmng
CGMBex8p9USuL0q03lwfVayhbwtYUPar1ljBjncOP7ZE/AYZX/YSvXo2GuXXc6TXh7AV7G5NXGZe
kAGl+9lPonK2zzWrpwXNlaEcxydMf+0fx9EJMc5BALY1NUhZXBwiKIn5CUf9TniIfBmC2LNvRAa+
1oTjQN1YQFjEXwdJJLe8Kqc+IEEWxEv0wRyZisbI0txB6s6MOxo2QB3fmZ5Qpk1XPnGcUno8b+bj
LexiQhpaCseCKq+y6j2u/54zF5MFQk/BmAGTaDMFjZvehizZgA55DvrSsw1tU/rd7+zz1z6+12+g
xXReg3f7JjBPn4nxUqqtP1CHo9d9c+wR/1YOwibzJcymoqQC/MvEVd3SWxrRdpkwUtcKDDAcNRze
Rek0ZM6rhWfwpMiloHd0aREhHeC0bRX/avNX5JFhCtaWkJ4qQM9+0yQjuRET5wiHZbaeMUb5a9mQ
iF8kQNdp9XMTK4X5Hi/v+qtMwkJXYa/yLiezdUq52eQF7p66ZMCxeVHIarD4IxPct8uuBFW9b4o8
M6OYhsOFmVcKec3zFrBtIK+IOcBsC3a235EZdl6cuY6VjGiE28VwjAyrSIwXL29HGPZRnnnEt/26
7f00qABSzdTVaH887tKoijMbwfYba3yLDc7Hy19ypANvoMHQ1rJX3tv6wwvpzjN7hfns9Rxo9U+3
X+k9WJp9vguCroDtDhidXco+M03vHT93X3cUY4tRHe8dcWzDElnsBjr0O7y+7uivwPQ1L4Vz6kup
tJ3YBaVZuWkgleyZzJNYWMSNAQpPKNZ/STTIHEHwr+GwN7h9pgcRFLzwPbRCJUVkJ2MMx5aBw/r2
cSXR/skxymHP9cW4j4Sp5OkHrcFLtvIKaE6PenH+oDAq2m5hxH1mAgC6gWEMsWuJiFo9ORxjEvdI
G0Q1uvmPb3KwjkCzB4mmOHOwPsF89CgnfRCO4jacOVbkKPF0d1jWyF4pYNDAkuvrpqr/VDHFKtjH
AG/OXZ++kEezmhwD7mZjWgva7jSzlUy1uB6HAEx/QJM6NwVBw8RhREPSOxTh7dlcTOglucmKQCcP
dYCwJ+yGC85FQXQv4/AoiTRt2GfB346erx3awzo6zGxACL+9VPQWTCn7AFnchh5PT9XwM9ZaqZdP
ZKd33LsCphWUXWz60BPRnkmFjVdO/9PY4xC3qRCuCgKQUMympNFu8MBMQhQk6iMsn3pqpzqVQffr
EjBr52WiZe2h/JYyJGDoBB4hVuI9WYy2qZkjvquab8JI/QuA8peDiSbpXW+H+SMNqvdyvL7sx6Jh
sj/eVfwvPgHSZSo3HZW1TvfY1X9E6FnLG/4D9Xv9V3dKWzCSFPI906OL3exA6Yaud2fzf8gLuGPf
Gnm14rb+72OmFIkPDSdV5hocWx10eOzT+iYycySe37rlxLv6NjF7aDmfzR1IYNkrpk6zm9VTyN2j
Y+mBOjhdZYJBd8uNPSI9PbSc0hJhaDHWlxvZOZ2TyUc2MD7A2pHNN5umD/u5B4P8YrYV+ei2lsLk
3c52yZQTDWahU6hAYYv/zjM79tOzSH+9bsgQGn8M8v2ncIhNDV2OKLscu0fH81vPwIATzTB1Ry93
+K0tcp4mBKPGTgggSv1eiVIzEtqA4kKc8OplxxQroKalOmsR1nrLMCutGRJKsVgWG+NKSl3urmrU
DVWTGTHpa3TD+QyZQhcz5MPFJdlKIuTgOjwquziPvYtE1LyMNtbPrdA3LooNEL6Vf3rjCE3frHvq
imVc8FVkpbdb16bkaRXyn72Pxg4/4WxeUYgB1T4JIOvDhzX9DyCZG0Md3mPynz81FbebNzjuboEO
ATACOvJs5oW2OS2/iSxbU9B4UtWd4TaV9WkGUO/OhH1RXL8/IkU0ihYdvzy89GG6oYk8t2wRoSrI
5FxvyfA3uqyp5A7LoUp2SEuYWbkFdO2X3jIFE8TGGFqvX69JEwujQSnODQP2CKvnsm8Jih8+DYLH
4UT+/Z+OZKfPQl0DKPp6wP/zYyQZccJU1R5fA+vYFrDzmnvwyjhBUp8taiJMZ7BSNvGp0tOlT9Gu
eOw/aTl4Ds9wwSZ8Ni1KpHP6HsIWT/iexAV6xEflLGCsDOiJod7ODgCuDw29A8ylDn0LXgfexO4d
eywFCevsA9WuohcbmiQQZHbeWG3q6ph1hYMSTr0C3psqDIAcVs1A2zrgUdiligdgcksTP/TGZW88
pyASlg5n7xMhWhxJjOiNuL5F3kmMeCjr3rHiemKnsMSj3YGbj86r0jc2nfKGdd90DsGTChv1N56N
W4By3vgF/vFz3jY+ZMeCv37tzkfFTD+LzsnVr8W0COxIr4OH14/RM3BfxgBz6pzA/JAr/8XTP/xO
yilekV5O7N31k9wXo03MJ+gEFNTBRTbOcNgn5yHlFBXQyU9aqLA/ftnO2V8DClIaz9m+GZkgNWfP
QPzQyId4zJn6E531AnOIgao3YtrvQX+7D+OjsNm/gZZt887C1TwM6hAtLiUtmw3VhKz1rtHhbVPb
J5ZkMlZwmUhAxDTAcOqkBN0WDxLjcCBAS4Aaf/RdRFxyLOpgCKOF17HHkqbirDcp3lt9lJxY64rT
ghG8u9L7WcyD99BoIEfURUH6v9ly/DQC/wt6HiAWl6HsLYyBcI/OjzEAN0qQtn8jjXkQGwcuk1zB
2EaJ4KSpEw49nuTMV+6Mh9d4s931axGfEfGD0RcA/+4rZGJWQjRAomDEY0RgbBT4yo20PJxgfGVP
1yEqhmjOQw2pHC8JqsS7g8H9pD2eSr12G7FBTo64JVTaxCDGY2p8fa9wcpVaQGXNxMIyQmnOhje+
q5VbciQxrIa+8U9WWa6fBsB+zRtjPwIYysHX+ghty/3Vlr4KJldHv9AutYuO4TPxU367uB5A0US9
rcSnY0OVfzV93fwfiRwolTNVgntzwrJfNcGaxMZXxMSzs7nC/wZxLGETKuR6jwWn0e5MmpnEB46W
6XsQv0Apb4FCPEkU9aylWjnD3Q4his1BpYc3PoJT/pRyh6kUfa+KECrJxpm/DRomFO3ijnJgEkd6
AHyYLfbej0Phet2III8gPzKvAcT06WwP4+tstzZdoYw9P3ucDsdaJTsCnxXpYpC8d4brwG5hc7k5
O5TnkefOyosT49+cyMISATY512M5qST8WEahwgOhXmpFj1wWnvAKf3xd8nf6rUIzH8kAkVZqtsx3
QTe4dVv4ZE/vakux9ADDeyszCtnwXeAYNsWFSs2dGQwieM3EugYRhu50Wk4yHikQP+f6JyoUsAbV
0fPLHnwhnSTXpwu77d/PGjRjxKnBqnvm4kc5nDAZ6GJhVXbgVMnycD8ZPWnUW/HHVBiqDY0VC/QZ
8iBdP14od3CH4Ja+yRSEWZMikZLNfDtlRXvTzFEyD2/LiRhMooZb2LT0gtz/tgMLlxWftzddD0jL
uXl5ugVzvTbwwIbCPp35AyJ4goYNh6CiOdNTcls/7NkaHOqrJQ8YGSMl+49dfrzMuUfoodFrvm/T
zkZkHtZ4UR1autkFwGsBpcJ3bqt1NdtpdeUDsPAcVoWVhdedB5/tA1y1UgAa43ADei6U/9S5YxyZ
yQwNkhjRw0boo70EdYP7dMYK7QG8VmwuNoU5cQFqLW3aGf9LFljqWuYG36fq3aKoNHDDh9MRN+fd
yQ3mbQz22vZpKYT+niYng0P6Ysyewd6p/eroDY8rhhnGacIjG6sXoz7WQ49bpWPBcVQZMSt2dkZu
ldnSNtM6hg3sl4Sj6W3cz6ZpEPlYUFDRUtF5wsw4tgISa3HtkxS72NQ3CfqzydtqzpMfsLWoj1pP
GBaQyBnc9EtuK9FUzO3fEuTitNX/rO5OsbpSSoDS5tBrBpTD9k4Q3Kf4ZNjRz0ykmlymxl+c/Cam
KFs8WRK3Vutv85nyOt0FNZG4finqrSfH9eC7wnxV34+6gwqI9Tq4TM8f7YbCNK7o6aQqVZJkBu80
c1VGQWdNLvLnJ3cPEcOqbET386R3hxudwESuQgPv+YaEj9KKc1VDp0cp5tKzWAl8ZN0EEuyb6bVZ
y0AB+Ys2HawbYhyNvTUbTRAmiIsgEtr7PCjmZmNSIFGY9WhmHXaC773UPhCW9Ml6EEQtBvygsICX
t931he7lMpVWxdh0aBAShUJJKHVpIG3NTIdZ+R1z6fogfULJG5YNWh5OorZQswuvwtqmUD7/NRhD
7ekg7A75G2rWjGSsTIunPjvQW95rRhqIia7lEQ1vZL6kmok3ZV6QzdWg3m5SIPXp2xAgY2DJOi73
j+BRjDwDp88W6r2xEZDpZ7h13Vn3LYL7UiCTfDA11Vjq/lRqmKDyTFg6T/d72LHjZtjbQ3OovIxy
ypyaZ4ESOrFB5ghKc9jUdvFfz/r93NZoS2aQ6if/4IHVTx4r3niPB93K+Q9MIzTazS1DrRztd2yx
LpdgrogwoaL/B10P7O1loEExAWk2V0r1uRLu5197CohXSFvP/eL4mVSv/Ej1jqeoBYPziAmkEBMp
v9+oM3ZBcsiospmkONCt0aHsfEtq7mnOSwQl/yNybaUwFzDDD526fV0xX0ruPz2gP2spCt3tRHtI
n0xLa7OVQf7HNwLpLVDko3f2krdOilkLFgsPUY3/LmmcGE2eCXebImn/UXXnyOHgCPYUwBpa2TGo
mPKXtlEHfylt9Eb62O+Toa3HLTvo8deXuYQ2Cr7s/mM9gNOkwCzf5W3KYne7oCL25GUeDMoBHd+l
+MojCfVvn4jxdUcyuIF9zQ01to9A2S26gMjiR4Eruxkh09A8FYEP/3QOPNYCs9feT16W+bGjvdJD
2PJRED950162HaFJavTnHfzqCJNHaF5pp9zsZQEmZH25iXRGveFBmxhX/zkIQE64U+Q0wWLlVIK8
jPqPPM27LTPjvwpM189H+CAofxQKJn4+VryhPRX7wWWlH7Pivp3Cv0h/fagQjH1nGZMXHO6c9cST
dcU1eyy5xvB7mQigjmuC440zq6OcG6tuHAr71rK2sClI0ah6rioVT+aiJJX30CyeZRzikDbk8ANc
NYtHqPkXp39x4DGH3lWkM5ZWL9SvtyAo29vcRYbnk2YuSgcHPHRAnjfQIun1Gjk1Qv7R7FY+g7/u
y9B5U1WXANC5NPVlthJDt58JQcYyXQmykrtkDgbG08jUgk5xPhiZwbbT5LaIqCbMSdS6fIvTPz/m
Uo2J2wTYKLQ8eWqRFi9YFwAxoHzULk/4bWPaddO+MZqt7NudSbw3kpq+840c4NGXWlNN+h2nujDm
EcuU1lpAFUXW7T5hPjcSO6lcBSRaJFAk4IqcutZS5u/1U6dg+zmPaBma6SlqjRLcbKWo4ZgRdXnP
+Lv1rEa9b08YaRtxt/vTzDECt+9HaXgAmqxNBI6SuRYimj9yG8DJkd8tj/ji5z9cI4KheYjmhBiZ
nhAjbym77ZMLbJRIWtpJzRGI5aND70ngdh1atJ17x+BXBPcEpiOppLhv2cZfxrGz3RAByyJAHETb
7f7bvCD123R26E/+rwumaghCV683YVAcFpoMJC23JKndePhYSkyncyMw1JhJWG+GplU6zM+4HJ8g
pWbMOpDGY1dkdwfQa9zfKZvweu4x1K47lAfabwheRjt8rhqMQxfQfBS6PHWhdTYuknezOEG9ZLWk
bPQ8npaZMoCuEkTVexaPqaHOkOvBnisg+ySJGrHRLoewVZyUOBJ4r9FZeQxXWpCi8dMwUkf3GyA3
HND4zr9ODJSLTd4XgvFEFWDltwvV/bn3pHwDhNW7ZwDIdorOFfohXzHNdPCj5D0FR+H8xZ6Rtu/W
Bnw5JuwEdNshQ39FgyKZ3uMCkHe77vl38Rj6Ho1GUMDrHTy3WBl3ApkNxV8l+MvVgh0ajdKwcx5n
mUsNMJ0A4Nqd7DJQ0jJqfNNNCzDONLMbTrI5/R5vjJHoDpB5+ynA1KlPSTwXG1neAQ5gqDgQjDir
wSNSoYzYuKU0em/puW1GYU2L/b5Sq86k+lO+CknSvcJhfPh+nAEV8GNlPy+vo5XXnd0v+dANoekL
SIzGKku0kSy2ktxBAumt5ceQUTyzHfweg5qYgz/DO2hnl/PyR8gyTAuBTWOt66iAsh/OyNAfYOBj
EcbbtF5i634W9zb2QMRfne6WdkRy7tUexd24/H++F3quPgYd3tHpaL35k/pNG0b4G1ejOYtvQ7xF
QEuaOqeLHThQ+MiwJ45ixHeCcPES3ZrT4ida+rSnsORTXdDnpmTr0Voi5troIxE8dp2JeYPImxXE
M7DtQLMNrorJJrdxr/iH3XNpzTm1YvZ5KuW2LJCZpSInAGXLHYtoulNycQgX8BXDvuw/i84ioZBq
ihNwImyNaWh5SUzIgKgWLbd5PrYLvJi70tnbrbtBwtu0j6ZUa4kDSIqZuzKnO9veKJ4wE4kgz1OL
PmBXF6VPxcSbSBfDCxOwTHRJDH3c9AdzbVutl99unUZtpDnF0l9NocDU6TnfL6FOT/RS3/tXnCfq
La+ZHC58INJw3T0BzGvbEJXBXze8LHGEydkWej8q/dyrArV4UYRJHh69T1jpx5QBxn7gb18fIDtn
tS2LzLN/5W5oBsePthAH3OYoBGSWuE/Q9n00m93SZu4xq7+AD/TUD8Kv3KfjjlBTRvqMsx99elxc
4Exd2ErIwODkJEAFEdGO41evY5Dkr4O0Lr3hnzgcrZojzSXKtjiLFJwVaWDOM2iZumSreQH1hRSb
l+ZJiQHxeibnKx3hdT+QRXhAufKF7SAeFpCzzYuU2hrYzcZerRZ93ESf37i0WMGOVET1RXOlOm93
8DDR76tcZQrGI75bYvqkR3WekKSS5bnHltY5W81kZd9/VADncMc8jnnG4O6W17MZsEfmdFGEP16T
1ZFn3afJdUW/feV1fmV0SqQKoMAqHAVb5vbKDFaeLg8OWgCy0Xf2BK+NXHZ8AlGAL09y8EeXS+OA
+6wl/pPQpaEIMG2aTn1p0tOTAKwEg3VVeBwNR2uSgnLbiEHfCYHiWzZOIxuBfZCJdv0D9Q0r3jfi
x1Ejx1nCHVC7W27nXJDm2CSHn95xCohafal1Y++yNZxsYf6T9J8naD+JCFE2VK2x78SNhdp9yhYV
snh2sF2qofROo9jxrqVuGXZzXJX175rogn9ZuoIz25ZrFGLXHhHab0Syn1LgFJ0KpsqNS81JAhWz
D225lpqpvucCae07Xg1rWaNgBO2cdcRSmXfntiA/GPPCLXNTwLiCOeDl/OXgyuLauxbCaUKK5XY9
3SFb0kXVDURYRO3nuTCzbM685obfD9/Eb8J1mZSyGT7ili2ha70SkvW0Da/TEQX4Sis+fbgUFJw3
6VBlU0vSPOoGiKJ54J+uyNaNQAIfSUnNltcY7G9cJUC1ZvoSdeF7dhvw/tLzRCpu70ErgHuTIq5g
1xjBzeAbw3owcPob2HOo7ZkGI461MknRLsfGSjqjK3hf3EO7bkClIjOb2yADt+le3V9MBBw+J3r5
kXyT2wENHy5y8Mr6f1n7GYko9pOo7ZbSBztpkk972H1aV3+oZyCPLgkCxtQZuhYJhvL5LusKKNK/
Kj2nAvJo8GjVUIGiwChwLoye4G1LlBEVdV2nO/yeX0wfEmmbUwNIbu+VIoYQarnJu4C+MgUofre5
e+zsXGKxKICR6OfbGXPXRSa6oYJ+dQWUZyAfpd6R0smPzJTlNUJDsumT44B8fLM0yx3QC4hh/YMt
TfhenTLUTKLRmU9RdVEW2sTcKBnYwsYB8LPQuEOgFI1ULUjeXOMQgrdxmzE5RWHLWSii99AO2l0a
Z54evrVDDjJ6QIEoU1KQolJVLOWGYAXZjO13EqBVctWn27jzbP5Jr7gfYAOUBid0uVSJRvsC4IGH
qu68BjLV5y9s+EdC31FOFoNv4KctOm6e3jV83/blj1y0TOd5ieMwvjxjd8/PiYLsMJaOexBGLo+q
vzITIfwtwHwhGSks2c15JJhrtmjxhQ/bOjREjfWkgDK8T9y3kRyY0rr+tcSaLahGurZjTz9XxVyY
Qtkd87N5fQGIyloiUU+bJFo1cyXWKhyGnUphC27qpRDbsLPYibiRmz53TlGr/HxFigPKN8uhv8x0
mTzSpoKLZ/4pRg03M6rR1Hlqh9L/05g2NGm83qKKFQA3+W+vOd4vySGpjZ3Z7R/tmZMZTnBiGwC7
evD22X/MCTc922FfgwBOB0A1Rj3d40lCqKHlv+MV3Ybp/wRB0gyrfp76ABErX3msrFWeP0JetFz0
KbwL8HNwcm+PvtaNvu8e1YqvwldcgctP4k5B9PwP1oBYmBetlk+277WF9zhsG4i11r10Anclm2EV
spy6VvBaZ6Ic5EnN1vJnmCgD/2TXdOQHRq5NKalRooWal8sbeDiYppIt6msNhNeHm4+av9u+j07N
XTU6vBRabpROwh6gLPEmEGj9KYSJ2yKKNv52yYocd5iASdLMg+1qTMcsC8VQ/Fw9w9U0ssn59VLL
FiXB/kebHoClU4jcE7llCMBW3rt5bbY5U6Q88IdiBh+67n/gDDv4cUL5udvOFCXqpN1Px4oyZD9Y
yD1QvKug8E31e4M99ve+barS5goK71gi9tH00N4qqksy1ypO5HO8/iQha4hEHycH2vPWDkiC9Hp2
e1+KpV2Aw/SfAypPx7kv3MvIYXyjNTTfpQ/jIL7Y2J09OGoK0pTZVqDsdN24x12ohyH06r6b/b1I
Q+raaR2bJX4rqVhlGAZmrqVIOoi4S9JAYPGAzb+ooLYgB7IKiQV9hWXeBLuXsqK0F8J1cUINR+wh
KU4MZ6/nbvmMpiXLEdTBwjdje+R59fcI63H83c61aHPPzRN7xr/mVJZ+aOu4uKn3wpijMfga2m53
2TIuKKRnqqJj3UFKhokSqiHrAjiUZi1fEmIuHHtJHKt3xLTTUDrOfSA42dbpSu7hUHjJqBIzJQL3
pV9JOEznW1GWs35QtoKtJ+sSDHoIYc6v/qw/7o2vyfZJo9kdIGYhC3s/2xXRWKvfYgVjZ9eDwWy5
6HoxiwZfhMuwfgowjcgnbue1VCsNwktegh1CHZvJkVstoD6h5KRSqUif0aM+M2Q/337x4ynXz0L6
4Ez/kQPcvGpLxiFUQPdUZ9u66lodY6CdDnsJeLrMBDJJy6r3+dkIgApwUsgsmGAIlv9Sn51neeaE
WTLRAubp5DItkQwT193ab4SmnE9/3sRyy+6tk88UzuqV78RZcvjIRZFKyqoFABlDukhleUpVUget
CGXlrAPSvviM6NK9uCa24s3ihPJbgULYB3a0T+4wVEi/6RyWl2qgwNtKhYlpLmI+eU/hYyMxuRwW
yngVz7yWH3iM3jACwCqrJ1KdvG09c17kl2Kry24sS0U8JLS3K6Vgwe5XLmLxASmAaTA0XnVr4PdD
Ln1IMcooK8cYKTehyN+M0bjYrqCmXrS3DZd7QpFmZL9+8f0hY90morjgacgViHaop0QTpRi14/G8
1ClciNScybN7yzRwBzkmLcXoC1EZlidjLkeQ9i7biS/wUpFHQePC12IYRaTkILaLJ8zSWHLwtmXb
meXNwZNXEW2oEKQGcxebXYn7Wf0q9E79IrQaHfiRkAWMdz9leNwKU7KkV0/v+1mCgLBZknYKUqiY
Jgzr0gL0FNrfR2+jdn7x3Kudhx3lAlQxwjgPWzWa5TVAakNP5t0rzvgEnIYQwqJa3PeY3hq0lZLa
3IObBpde4FTq+MVNiBYWw4t6rZZDY0TFEHO1SYWGRLxRRygvGe/TpAJiz5g9KJY06Ib0+41uT/JC
6+dbW3LMckjkl2NM/0ymmQ2CEUdUoe/ZJLJUIxTntnrwXP35JjJgeDXQhV/Nqto848H+3cGEWRLu
2R2+E8aL5n9KaXyBF/rCgPfdQqgMKdO9CeeaZnO/S8lDir8kyfdyMxfbv/Sp3XshdsK/l02kBt9g
Z1h267yuhaK+BzljMbvTJoos0qcuFF/lDY37JVRgtRMQd8c3CByNX2seD0aI1NZ7LksV61QXumXF
TOOKXThxAJCR0SZddG5Ke5KQwhKZXGUJq3VBQ1KOY1c5BNFtXJunH821d8n21wBssU3zc7lFZlhV
gaICOFzdpngN6Uw4lTfbuNsUJYVX3V/wkJkWbo5/IP4pO0hJyl4euGE+Wm7xe0c6zaMa5NLB1s4s
cqt/vuOK9YDqHg/DwFyurZ5MQBg8lPzH+Sofa8YjRSrP/HjWMAxl4HslUpB63Yz8+K1ZnR/uryMR
lgN7phW8bRziGcdDA2bQ+whsiT+PKNPxK4HyrVW2J6mfRdiG2Yywe6poUeUFH2K+aLItXWZeD5uJ
XzcyNIvvFC65DAhIX1rZOquWLfZFoHjR15hYJMkruMVkkmGMv9bOA0vM47x7yFTGc9ZmJHh65bBz
QYJQh3y8xZWpR9pFxFmN7YzUYEGbk+O3yDsUyGvseZDO3yhqTAMuJGygJaAC0i6g8CYeoxAgm5am
WA5jaEazR2WdGQzIO6+Fl1LE9Ry2aMrmWLeg8UL0kbXSvQyD/5Y2uHgqWL9p0giyza1r6f2gdjQL
uRr8Kgf1wysVmIAXZ37og1uyTUexbNdK+dNNZFboOJkBGDYz7rcKw6Q+K9NZOufbgFURD1ZrAgjn
dwrzAbK0O48c0Gs21NbB4hDeovd9GMRtCmrYe8ILuGt7CTX5yDyCYM8w55jGvWSerfrTLlL9M8WE
SkXujXdRp5Pv11gWVPgVTz7IE6fhDXI8Obbzb6MmKLA238QLcwdtiADVbrVknR4fQWhRs6iglRRG
yXzep6h0cCiCXQ8RlJKrdcuO6tevgV+prJfjbKOlLOnh9up8GXMatDTW13FdknYFy6nczFSX8yny
YbtVBy51I3r8hUyvEgO5O5jWDP1Yt/P3EIZWt/E0Fa6X1nXdO8ZejA2pDA1n0XzlRIX0/HLEzCdh
ULr27Ew00SaJ8x0KHUxKDKbfSBGKz2K+oTuLNxWHyBA6KpN4Wz/3MgEA9SwMn6KCypyk7xzYMEj7
cJ3kwNzDLKyyp7bszqKr/8bt1N5/McfzLDU46PS/53/VcRKYuIkT6pahhn4wqb+ZuHHvrm9OohFU
ObXEugkqZtWJDuTNaBCuL95zP0JdQ5ZctmZ3CicA2InR/yrN1iCTQ4OSoRXY0X3JgLqnWbsjpBjY
OhsT2p01oSoKafeDTib1GtY/ra2oOrRZdLdXVz2BeRbv/z+2sQfuv8Vs2RXvhQ0n90R3v6ojrtaW
DBKChx6zsfG04rGoXPxUsXbbkiUNeKYaO/VkLeXodB73GeWETiCr9y3cwuv2sK2GvGm4T1dJp5hy
9A+DdY7Ot/ry0K1eDMWTyRbpCKacpEI4X2lRt+Oyae2QF+qb8O0P5Y7FuMWs5nJiEvSZC6UEpuSQ
x8V6FFzIHvxqSB9fiVW9rISIQ+bxghnuUJHra9Pyay88MQhft9rRJmcAqRZIKcyKrCVE1tAef2do
VVu72n5/m+wWcCXEwOsE+gPNJhBMyIz1OV7Ynk1aCvD4WM2Yh635RdJaHv9dDYWZ4G04vskyjmKT
vzyEbMuXYz99HZiiPIrfxEkw+RsMOkiRmRywnpdVub/6LQ+SKLRLpjQYpLz1FC5C3OWmnypnM9cv
zoPpuHxBpsKBCCMOSY+6sso0X9ZwJfUhDEtK+er21NNYuFMGRx0nEeY5Vv+gBU7oyelxDmxpcFRL
ygjbBmx18P4mz+EoE8sguKLG+Pu4E041xLWCbLvaN/j66yeUOW16/cAO3RUwRxor7G1WafdGd6Y6
PmbFGyN/6bhD5zPDchrGLLITy00DkAjLEvyZ5gLDk0xFjeyqVvh5nPu8J+REcADDbVXKcFHs/ji9
vsSAJQb8SM1L5VYnyVu6m9+v349wlrNiCXqdZ0l4Hf9Df2SMK+gLNAwbXWOoeei8eMFlByFe/pX5
QYd5jjBY90qmJFHXfUVONg1mc0osUOwNC6o6FiiSZuN6DCtPyjfVFdgQ0zYJrZEft4Bwx5z8NNVw
rqZ7uzfHdVhDaoraDE3OgUEIIOWWafVNqYQB8jU7cHJeYUy/z47Fn0SzyD97yBiT6gWCbQyOOk7E
dVERAlB5ikiHfC711/yTKk1NpFcxkOp2jNTW03VMAxirah71eC5pldTJx8UCZ1lULz6VCQkTq3o5
cgmZqhIE0zNTv3AVankAeCFuTxT/Fg+qGFxPjPZy25GO17fBRWoTNsxN8bI8hhVdbIPPn2qE8SNb
h6lmYrfxCTVC+SzdjZg8aCr6roFTKZI2oSyfM327808Dh0XoD95gqXJxCCXXl3p3YbRCFbDzw43F
i4arv6FjXOxtML8vVEU2NjeH277oNeHvi4aNC7DS0nM67sb5opPKCZwh3VMmJY5PiBlqh578+vDX
D1C5ZLGRxOLnw7U7SD2m7u04qRRaWNkcZQcfBVIZu6Szax4zgOYgBjGTr2GdmNeUY3Ti1wjO/Xhx
iMQS00IFFvdnob41FBa/R6cPKWZeOVPmZ2oBfKKmlNSWZWKUYXCIKJ1WHCd28DFwmhKfhTUDgUwT
nruKddzh5F32i5X1LFetkqKFgTBTPcLkvWh2qi/0ptYgfSjdp3eNuEId8C7Pn4C99vJN92VWPtBF
ToabB0DbywDC7jf78LmdwvYOO1D5UdsGxvHhldlE8gM911Wvv+JMs+dGGT/HHDmNJLeoArnjbFTy
+hUF2b7kpAcYxL0V6hyi0XtKxVsIwO5homhLUQyV8hpfkQFI2XndKWf1u/pbfIJ82pNdJuU33l/7
MeMVo1lrqX9jJlqUd/h2Y6+nX/6aWo6ukzXuGv54fV2/JY+Byd/Bzz5RchpZlasRz/2zq5od65gN
mf36+EKQpl5nm+km9Z3Z5TAt/u+eiPQrVejG8bvKq2ca2UXp0Zb1CVjtmEMZpsHiSs5XiLcYTLBP
2KLRXmJY6nN8JTm3mUryNGay/1qodTcp33WeXiKOmvai7c6vJ/sWtFrjSHxgJewXGi3XYSLjhplM
f+wR1Gsaf8Hu/CNCDSbkKxfDTLxlSSu1XHTqKb+e01XdLvfNANsOIIALiAkbVco8OaLG96X7OKAr
zzIUdEvdqxups7GMNnji0relmo75dR8XrFDM27J1djfqrgxio26vyFBOlgtrJPbVWQTxjtzdYSTr
KTdN6L53gRMX7MI22RL0xlXYErMZfF40987t4Bqc5nRxUzTtFvvN376wHzlRZ1FbXVsZnS6Q1P8S
XEfH4UV1F0zomAo6AwNkxN45zIbiMUrA0dcqv8yU4+3WQQ9kwaQxM8JpxewClAbGfOHIxLFFO3oQ
ZRo5aEqoCc4XUAYcadaeBWbI2KOzcpjjwoL5c4yWwrk9vRoKRxcH9Dc/ujGPEXD7i6/Z98BTDNBY
XVHY8NC8JYvnlWHzQsenZw/jpO4QZzOwTtZZVNt/5FOXQgCLYhn0ftfA6OJiLmJMXAkB+2Y9U5zj
ZzGkq6vQU5HJ4nvsYSsRNHTjbyp6IotxoHBAUW3BYLP0O/+8smsRKqddyzC0fmhGf4I6hEBgwxqU
5SfBKKoW5pDJTSiU2p/cA0IojkJp0X7193RchVnDjcc2mOzhKPTxF3Bgr3E5Xj0L20Y5UsO9fcm5
PTEtZVgl6UrQCKyj74DXB/BnDziCFPFWQfLorlnIWdv0D1HQp3+pGHgJCuLzv0z+WodMNCNM63zd
Etp5yv/g1UGr/Dh+zMHETBb0CIuZjdYysc6yRzSId0qoQIp7BR5lrUeS6y89cVsAaGOaB7/emD6A
MdA2+t1oJ7dR06Imz9cobEMF3940QGcVE6H7h6Vx1sv2DLN8GD4huLeTrVgBSoCvqlghwb2g0XoR
UPgOhb4DMKm+V8SJT4ByvWkr3fL1A8YkjHRb0dJKheGHqJZUf7AkYKHZI+cgnjMYPIiJTBpod+gd
xXxAw2D1G2YlWLdJDI/mZhsRrIocEKxTZKyrG5yfOCaHAsS+ZFEEWk8rzzin7koKS0j0+R7YGsxV
AdbhS/3FaDvMB4OWLzzUbtKNN7oB/Tpn6gTV3c89z0aRAz4BAjBa/kJ6zKf8/V9zMrmYr0ZoDbUw
vF5WimPSEzZx3kO8q9ukAKa/WbUzg8JQ/Fwc0pjFXGlAR3xnErYyy8eMb25kV6eqbYfA2YQkJi6d
reWZxSqiP9iDYOU8M0+RP9ez3HkWSrVacKH4G8WXLY8l249qpEUjhGY5NNaEYFOu9LAFUR4kkiAL
e4kyq8jt/gaPk8uKkA70Y6YpwzF3aW7jNZ2DtzOl7ScLPx1E3HjwjeK3JW7QUVbony9kOLphtVCU
fwfmjretNFrkEpT41Wqky6NC8YQAleTtEbFFd3kP97NFEasDRG4PLCXwPQMb2NA3/ZoFGJlrXHRn
6I8VpcGKQPHAKg3wcOaRIMV0FZUKquM5kQwXJZGklCiDk73z4pOCzve7CzEm8iN3vcK9uxRujsmd
8tlxUmArd95uOn7Q5fu9RjT5jCsVmwdrMf/YyKyqHlHs3ytmDRrnKdVqQTAAAht9dXeORbDZrWYs
C9r85+YtfFFmG5V5QiC0JEW7DLELmV5fUhCWxQQIxTO9+YKwi+Ommp+wHnh9ppMUGx7wcTNvH/Hh
qaUyWi1ONy/KpM5Pr0ZndCYtf2rVXSMJ/iWkefPqbdNsY5udEFXm6/eAduNgDVs7Hvm1Q8f//NVf
o4kS3J9lSJjzIAu/Nya2OhNQMZ1wZon2JdkEOPddo4yI3RQtjseVgGpNlVrnO8uj2jWzwxiH7uzd
FRAAiG7Rl4NQV89UkXUx/CUPznw6NHf5ntCrCUAGsxMvCugMjWCa6yldF0p06OdsnrpvIAQbiRBl
wVa+kuJpIKIRhR7yDh/BAiLPSpK4wyRExM7jz7521IYueqy7zhOglznfBds0g8b3iSrspOnC5lFS
M4+YqLrD6ZmcXXzXoC71nrx2OwtzHoZmCAFR0EY7Ze3QOKXF9TF7ocrLMtbR7/FpRPyUUehFrjg0
IXD3RBl5U4NVW0YaHW6pmteG0qTBeA7hfhIpn/UxHLE5cmY7vi4BL7d4C+2N4c7CoPtbd0Dc1WvH
yUzl87OG45aIbm6D3r5Cr3qXqiMODBpz9ByXOmS6oy8EhaokAbzbd6QmT2T2iEW+Dcpcs7eeERVL
MgKu9ixXra6S/wcugNTHxdqq667piFRq9cGZ9DyDP9WxbsguFJ2aHOcV0DXanKXFY4HEKVzuDmiY
Dx06jJNvtN1lVgBTRnPwvgEyGrO8CM7XcaQNnr+XHwNVa4mMfO5iOqa1N19fFeOuKg/6byWb/OoM
94dkFf/458BUQE97lSLhp/eCIxCz9KDINCe2nGsq30eQnPTUmOmBcrmJnTqbKMgLtO680FDaa8c0
YjTIhbU/p+igD2yPlbIJ5EAIcudEihiTQKDtnq+VEdJV1Hz1zIzb751TBKoueBW1mm04hmkbiNpw
iGZq0MH+Rn9uMPKfGtljLZyBeLnKQncm4VUTjuLa4PCxWrr9kFdZp/oRUkwTa/c/xae0xZx//09X
nDTbzADdMDzMYAVhwhtqPN3MfDAufuaxPTHapvvctefMyKmv6ZFQweNPHwOH/acs2bkxaI9V7Dfn
NP/763xZ7eTQRoO8wuICc9/KpZizwOaWLGzcxKJfE4/FAvLnRBeI6Qfu1xsbOCO/n3tg9cbcBRDY
HQLONnygVJ34G8wcnWe1W1F9udJrQWH3vtmZ3dSTqfPoV9HhPk4QuznytdnO92++85U/Kvx93aBn
uw7XiPxJRiXziXx1TvdR4SxrkaBMkXE8+UTj0wJKS5GwJrtDmp+DZkVyIXs26ZA20/KdCA01p0gY
T4GFCNGjl86PrS1j3B/XKTzzapRceFbSoJIj8Z/ardYDKINZdQ0cVTy2VZ+ufVHEyO9ZbMV0JP8r
qCX5bk8BiS2dpPA7k4P9AcSQtAEpL/RqYWVxmRbsXEvJ0w/QbV4WTJ3SAxTH9QuUjP/UsCeKIxGl
5A9Xk+kRTMHCwItdQr1o8e6n0pcdsEmgb4bs1qW6kgX0CpJz4yGWeae3vQQJDEjHVVu5tfCboDHa
eV9FAQGlkefT4CL0VSviP10CB3uDMi/AJBOenNru8GnEErDjBbMWl+gR3DHyELsuFJDU4f8xKdnk
c1R+5soNx5tmgpm95Thgzam+uOqE2363eBmA9puS/ubYqMiVyHFODH18QaoMqYHsEfE9UgkBPy7Y
y5LbFi7Di7R6RfrN+kUob4/vk+sqkFNd0s+sSvhfGZxU76TT67PS+1yWJB3J8mhsmFLFle36Z+Ba
qFL0uR/fI8h/CUuiYcAEX/SaW9ME8CLGyukzBFKD9E632RN9VMAsPl7OUE2lx9fa0fMLQ+bx1RYm
kywaTz75v4JGHWG814wjVNcHpcfjZRQ5++4mQw2rm/ZvrZmz4QwOaNHwjp/QsLmqBF9Go+2m3YmG
NAgZCNQ6iiHwt0XqaU9lQuLYTByTmCOqe16yfBam/i9sTOFkOP/Yi1bsJCCsIMmP02Vjp/YPbpSb
ua5krRHmEeL+pURsEn69Ekn3fLo7m0aEhCFUmFP/hHKjgz2c/6BoXuJOsC4tMO+Oi7EEHIxpMPmX
z8eWmrxROgvIGDqI5wQvU/qRJTRrVlbGDLIPGlTma/haWN9xMegHBS2EjU7YgnAiyLju5AubRTGs
Pyl5d6L+TcQQh/SYjQ5LaYtsUo5aLsGlupMrvQB4koRv22b1siVBFmMqnVJS3Ix+PLbutth+yJNi
LvSWsN+w4hIcFAz6/nolBi57BIIQ1sCgHn5Imo9Jz7mAznQiZN8R64SXnc3ecIlKLhU+tt4Pm9wc
HdgHYocgaumDOaVCFs+k4QidVGUHSp2kcY+Yu9luCUlSBzgPBpqnubMiLXE1hfUN4nIxDdKeXFAO
t+bYivVNBwtOU4FhncYQ+SgoptQMBZkDGwD90os6KF1SH45bf5uUULqiP8Q8ztGmQ3fRsZdLYvaO
0k5S+YovFwTsaQcJSA36B/HrcgY5R7sqdYB32AKqJmMIkgYjt/CzRsQZtF9j32tR01VjQXTntLQ4
4zG7VP3py0Ua/Yp/nfoIj/50iGMgeIS7HsphwGpLIJ6rwkeNMND3i3PqNzAPZji6mW2yuUqlNVe6
6fYPTrhaiqfGueXDffFVEsFDDHQpXjSlZT38eK8WpamEiWL0zrKwaa2pBZsvX6r6nHT5UvMP36Df
6L+JEO0BuwSQEMr/ZMgM85YoWNMQMZ1RJa2LUzPHgn5Ihw8Olp0W2dsh1nKOGzS3TUvoYJ19Z15a
5GrXxeuTKfPuAulYq1EE2L2UFwS1vWvZTvcJId8GIc8b9T9XXZthceEwSX6Wny0B5n3GsRXGmhlo
G5jVev4kdWB4cBXdtjlj4viCRkPnw1k9UQskGUL1yJ9tVfZyBegY9aFxvjIW3wbFHWvOLprJo/4D
HyDO9/ymU0gzVptJbnguiuSLW1JOgp1nLZjR+e1CCzA0gdl3fGk355SW/nbp1yKnPqp6tTLdJG/9
FY74rZMytfjGAPDt4L6bsDAXhbMlZ9Wo5i7YrrC4SPWRGfI6sDTfZ2/Vtrl0hc7JwPGSknjVqS/4
MD8ehyz47r0pklhKTYFsglu+dj1cHlDo7UYsIkoYdn0o9LAPstw7Me4oirCGuTzpjRiN+1xT6Yd2
omMexmbnzJFS5D0CwzOVbHyUuZD+Lu6Mr8wbBj30lb9Az+Z9ak4F21SG5nAsIGlxZxpMU7AodUvY
+lIcf1Q8YB3scMzqJZGfTguh78V7F7ABqNYcG59YDRwOkpuaOmzjtUg//bplWanuaWBdavQC2PCj
Jzs+CkAMOIP4j1nC8ro4/4Fm9LX6fOlLuWcqJ2/LKWohU1/1SV1pNR5mBTj332nnyi7rUByKdmj/
PXr+jizq/oupqqcoVKnWe418TrOa6Q7fsynFaxuLnWp9aqnOcsBS4nC/4QCaQeP777x2Qf16O51N
0cRgyYyGeDmsHWVps3Ows0YwixX/QkZoYLoBOT+BQRUdf7PcfP07/Qph7QraDw7jrYISMWHQB4P8
OxiC1bJzFyepQB4zFRlP2vT78E8w7irWxSq3DfEuPjWLK74j2eiIvsrk8X87e8lbu2Gio1Tw04+l
TahaEM4g6SUOhx9pr9lk+4AFh90vaJqNJYDpLyXhHVsnvSy593MD1I48bUywVBpr3ZeB0qn91W1N
JQY7NqixUPkuUCGlItZgxrv8lEFSDnwZ9qRnlaOOZYmdrxU7DEvQjYjYnrE7QcUevApKSV+gjEOH
++Gg60CFCfoiD9I0TtguYFz2z9marJfVYsmTjumzS7S9xMrAzPQjwws841R8PWPs/qb1XTWBCBfP
kUdU592tVMXgudY7eAhVCB8Kn/87wYLtdOoxr00F356t2ixUrnKHZZVlc52NhPbfWuiFDNyIb8fo
Qd2aXy+0b1NT7AmFiITSulGTtadQ8Vasb+oKUJsf8So1xdZDr7WfWetOC3VlbbdriPWITZCRI1O0
KtlwRU74XfPPhbiNkuOhAK/iFS7IYjUlOZfTnIrm6qFHONSv0V6sHPMsZcLIoulscvBQ7uynp3bm
YUzNsVrMN+E+sSNg99fwX9o9YxAvodEqLyIXNTai1rhX0VxZowA9jb9+sx3Bd4MdchHV3LW3n43j
uZuQJU3uwCV3cggR6Ki/Tj4VDW+cAx1QW+fYHHgdOVSWv9UP+tKrgKziFUAaaq4ecxv+9XtUOJ5n
cd+8fdmV0R2s7vNcvwAHPjPFpl9+Ek8FLg2xWO2auWSoOiIGvxbEJrnjUj6+7DwYIGOCIhoiX3lR
YX12hhaHugEOgEIwydOhXHg8moT98b4K6s6i5Ah91QXKDzlM2VtN2AxwEaiTY8u4LPkJ95Gg64lm
4CNsjgTrPVa7y3rf3kZeqAGbOchew4jXkWyxRA7Up3Rg50UFwalYWcKpQfeIrrKXmHuVbnsj+hmt
tq2mr2zvCioXqwzgF8jZakfuLRo6kkykh1OWY5ZakCMpf8kNH2LTTIx2ONRjuTn5Hfl9t7ZoveJv
2acc0y7xIfWeHS1i69y9SlgXcx6ZsapPlqGfrFsK80M7CAT34x7npDuezZUs0W7ApvAp8a/wPWch
JEt/p6SvKuItQU3tJRF26C/ANctUs1zroSg2wDcyMpfi1wEvJsny2XZ29sHzDMNR7+MLQZUtExPn
JS2OJw0i94zVcn0BG14Syhfz5NcnSt29d8yfsaDDucd8/ES8TdOUY8Ss62E44GYwjoYv+iRU3auh
XzF4QGGinOo4OFA3ZCtWLfutbGMwCJnSEvMHVg1CJ4M0jmGWQ0Q7StffVlg2VmhTADvU9DcIeU19
1XQ/1bKDRv8uEUaVtWmKzsVoua85FP8OLi9tgobNKLFxK1MCzRD74p5O4gE3RbjZzhp5U0jKwQXP
cOyU502LxzpzPERvgUxohlRFUEOcpPkl++Fu8/W0WOEP7sx1k0+YOYDlKnTN+MGgGd0TGols14X7
1tBfytlMb5ma6jHhG0M2nfeGvoSZT1qIcKSSPw+V+yO1u+c17jVMlokkfgfZ8f1O/0jKtUI4HsWk
xn4oEv2rFnmBv+kS8gePeq5OtaFk9Ns54QPtj1oVQLXFJZIDGDSxtFJB2J4AL6Hu5OFXbj5DCiob
UhaciYW32R/Ri3J7+u++iOMe0DdrA4kzn0lza8U96ucm7SzbLiLKWFb2vUUEa41/1/MGWp94cJGc
AE5nnEelw9aAMmcPUPh7CZMYjE6An7N/O2DQPKaE5rUSzf7qTqS5zYqjCA75TR3x3cLam6dV/nOz
KnlqdPb2sZCuMjH/+o+gAMYA1lfCAjV56aV3fjUhjMp3ULEbNqaXcy/zZJcLulF/OVxrJNrx7qJK
yaEjD4DIIYUC+To8F3jysN9OuQJ/oW1w1F6iqfWkNF1a4jW7QVNgPi0qusKhZaFxMHJGRiR5aEkJ
Fh3XLy9PFXbe1JvZyusVBgf7YsbX8+8bc12ZBtiGXNkoNaFnEaa6DJhHi0r7hUqxTqASqDhSTkJ9
KWS99JF1xcvrfxTuH7DxiFg0KmOx9AxQEM0GkiVrRp+kvkdxftiSRrU/WXCdUKitMpTkv9McvC6Q
GnEaza2my+RsmRgothdrKZtX4m0LVdSdZMDI229+PuDovaP+00FJLhAwET0LUaXwY0H9ZMUiuI0B
HHJ0ZwYy+MEhD8GwYZcpy6cs/fdzS6NNv4xLQPOPJ7NUERi9Qq0LOA/IGaQJWC5J9/HuvFlpz3yW
vXR8gY+3EipYGSKOZIoeWYuOaTYSRTf9NC6oEaTH1WmxzYYtmdZACEDM7N+bZtCSug0I3pctzy8M
VMCjK0jFg4eUqUD4Fj3KinINtrQYHnSSQfmuWalOg1G2+mZ87sBNIVhnNfT+4yj05orSMqme/wNF
JViAKr6gHRrg9Ch45nJ17g78C1vmyMF4vcXm5+YREq1tL45EDgjGSzo6axsPgjp4YPIHO03l8tLH
LIaARvfmV8IRDNHiNxJiUpvzjyXEXzpWSJ+6zh+3Ut2kbhXYCHo+F+QULo+1VrvyX9gGVcIqY7Od
6GNi629eAA7bkOMJCPw0dVWffiGLnoG6+nI7w2oAX8NVtE8ONhSRu72LPVXZPQwFMJ4/aDNcbKdp
7NtB9T8oXMig7E83QWEsWbfLVw6lBClNbMYHBeebnt5UMZsTP/zO0r5EPM9xvmGV1x/HJHMLPA1V
pggHeHmG0DqHp/Uncb7ona/xQt4tYv3nNqqoS2H28OlLkCSybTZ3oE+Dp9Z33PKDlFZG+A2uu2s8
G9epkNtmMXfoS6Qt9kAivh6fN75yoDAg2hxoAX57LrIYQ1ZYjshzaF0S9cO/o2bmtq43LtCh4xlq
5i3TJFDFyyl7pOy/DkeqfuZGY9bqkEZwi8aMmJwa89JglZsip3EFlgcruiOY3rOE+XRXfH3rCqxO
NOuG4XK8RmjRQv2vwlApUXN7hFV/e9S3TIKs9U53QX6przyjEYlTaWmENyF7LfxQn21aR8mnBY3g
QlLdbj22hwe6gcETmcBPVIEAxN1H2TtARgrucwHBLOjDAHrSaQRWZwr+80Z8V2oejGQb5dOlFLRI
sy1TdSaxBJuT6JBeSSVh32XmWMG/KsRsEbXcGxY8p58Nm7eiw3e73wLq7a6gywfkow5gMuhYR5kq
CHZoutCCCep1kr6Nv6czBr85+UIDwb5Q9n/N5i+MYmqtaRCxgpgfuz0b0rfb8V8X5/HlJQLQahGv
X5B6GNvOzRo6oopkMeaJIXL9SCTNPRtX/wwKv8+HfKR1uE23bJ4uCVu5F0zf0h2OwWO06NKDXLAe
Uyk+Wmv2pWwnZOcELYmMNfG2L9i3WDMhxjNb/d0wdOcHubtznzC6bRemj4kFTTe+10fTjTvKGWgw
SuO7p5JGzLAOMRSnqYoDRnOdhKfx8AraXGNKgeQL9H5v3VKhOl4JLezWg6OP718CPaSpXcrhOSuX
KrSU5k1Fpr/1oFRTjPj77P1BKEHN/Rt0dP3bzaN85K1MxrxawnGcvxJkGkjEsiTl/wuy+3VoevKH
+uC2IvyuGNi1VU+B39PO8dS7ohzf6hNgK3Yj5eWPPbUlBY9Gv788xT8Mug28/mJl2Mj6cN0bgngZ
v5W6u9TntnD5+Svw2oSlLfvHNnzQTWgjDwCqo2aK9Lx5blPsCUFr8V0BYewucZHgGdY/P61Iz27w
gkSt29VevyvlFVhg1KgjIYwCnEIBvsZlenSvdwwHyVUGRVMt2wIOmU+9We96g6n04sRrHTOpD88b
5Wj+lcXYnTVDv7sz/rfiKdxPNcwehGcjHNW9fgG1zBGzBnbwTbceZXdTM55xsI/H8m/mXufxRhQz
xAcK/nOJNNjsoupgf3giq+Ifut+noSV1U0U7m3Kd5Ut/UbhY8WxUUm2ExesYwpc21Iygj9beeIve
Jgqkv23oLE1y51e7bFvc+vmo/zLA7r6HlxzkLyxr8xPHnaw5sC4LSm/JORglTEO/034J+geiVWa3
nX/c4bUu+CErGVW2mLZnnoOk9XdNIkNUmiQRyWplkdZryQaut/IjGtInyCqpqQlYLKYmv9RCDGpH
whF9nzjrCFDbClPjK3kLddjIgGFsf8D0BhKwZ4l7Uhf25pSUkhOkLbTGn6Q0cwKPz0wH1zm8o7t2
t+O7tjENTqaIZpEVpR52ftZFW/TALIn94mXfgRuMig7/KA9B/UHgRM6K0+S0J11vZpiEhjFlCx2T
nDbsz2HJc/y+Zrr7gElcWB3KOV+jFTnBZeX3e0mAf8x+W7h737KdHbuUbo7m/6WjEVXKaSqotfra
XsalWYkT0OX0d5FnxLZp1C2PiGvS9PsDQc/oqXEo1f+SROeB3x1ajV+TPBdG1qnBrPxcslehS5m1
4/4kE/fRCETk49KNWJ1hswc4RuUpd4G5oQtUzjImiE+fRSp7HcPVJiu40be7UfReXNcrCou60TGX
YoWsh0oIeINZDvi+mBU9PnEHsBzLXxnNP95yzqN5zBJTDE7oh/wnITKhcTq/+hUofTq3bQAk+/25
Jnmd9YxJLtG7BKKviUVs8TJbFEcgxna0xy5Tk5ycykLjM/onZ9y7TxKO/nONbCQZuL/W6g+ZwyjE
swM2ZzE6ew66EpIZhIJAuAbnESMVQaY2UDu1kpTun6SMt622YE1rnHWFZxg7BucRDTNGl/lgeUfc
drHwLa17O6hU0zYZn5u7Q3Bwhdvp5OkBi1vkvOZ6QDsPhCoChnNqjx9y+kPpyhAnY/lf3Wem4OiB
7Kx/5fP4o6f5Tnef+oHA3ijCSnq4CN38/lsmvpZK3Gj/CWlEOic9cpZBovaCd7p0kZypSEV2Wpf5
caqmkdWtZmwuvppE71lfUdRLt4cbz26Mm6eMucrNRp9dMLHa+rRWByYlCA11XAJ6jvWPo0gljBHh
51XiBgGsW1iZpcpS4UsLn17iHB8CzdIukWVdY13wwqTAKVhWLGk4BiCmuTbMSFPjAw1ZH6KXF90m
oQT5Iz390EZLpn0ZdkiS0dOQTlvK0fTys1WxDKdMR5LaBK2pn+aMvfiGqDN5PhhV0SE6Cwqqe83h
3npSyyMJtHQEtOBV+jLszVlt6wjOvGQrKUad02ChlxYkF900PVFDoMDukH92N2O4foXUB67FtRu/
+PmoW9xonghM1OvE9toVv+lLQk9JVUUbcJV0u/wlOGuE5WvG5w9q4c3BtokLc20lumaYYXDoyfzT
vKyjtmHHYbCzwPTGh1IyquvviyBDtFgogXLg7B+WnGWPmOjt5TQHb6iegtBxLa5oEyrTBX8yHLCB
FWW9H70GkZCS4/XIrmtAXQ+4zpyUXnjELidfwdyCQTQk2zf1PKdHlArR10dEQXxXY4+IJUWkJUUv
S0hIimiLq4RXBg51Oa1Yd3BNhVBJvQBNVJtmEmWb8feZ/lOb48a2T+SQN66XTUes5hWSp0oOlRiO
qjfbU+4zmVNZ2Wap0L5RQFCP+RnQo9tH+qIk+GscXQabW3hmBTtHJJKlr8BMiriK+Qszq4Kn8brL
0oqb+FC3ix8CEy2LqjjpexdJPQ+KIz9Tzh/sMr3COSNTDV0mTE4pClmOSlERKx10pV/3PgvbJiZW
fZZnKtfh/Q/kF0Ghq4ES7/77TTarJrh1OUKFbHZpYiGwd3EdFCkIvk/VzvfsoaTFbBKD5srJt0m6
taVLTQcPpI5wm+jqEU2hLEqqWPMhJw+eJAgsIXInJiO9/aAW2jJp4zOkqO8kB7I912tFR1KvHn2i
A5AID0uViIbTySlCfoLEgFUwU/VFDjD3I/SDv36o6xvlaocKQ3PcouSLB+kvPZDO1Sweqn/ZVUcC
0l/ME+ewwUrgLtJ3zUO0f2Nemg1j8wET/oY6ONOGEZlfyC2A/deMIqcdi73hQXbEFsUNquzy5jdY
R2819CpTb24QDYeZjOwNz4x4znCtekPW+2NFhZT9nIE536l4m4IOHmDezSE8aJIjcO7d3FTrsSxC
kKVNIQd5AuLALzDuA/rpN2m5G1e70vCmuuGS9rf7ED4iOD0Q7a/EL4/HynNRA6IXqhB+PJGL26qm
Czvbb6h/a7vK4SgjBYkuwHjthUOn/mW2iVmyGoiOygWnX7IaLdluqan3L8Z6rSyPysHsv5nkrhm7
k+Y4MtE62LsLck5vrXGS1SQ/4fGpEqK0X/VTXfb4U5GCWkd4jBetOXEAqvzFi/XXheqYX1xoV3fh
dEeRWIWoCxCfaQMUlNzne1qT4nNCnEvN8y1a5Kq7qSWhD/BC8DInMkXz9WQXNlJuJixBqKp8m4B5
CsZ0QY77lRhhnqnrHDeL1UksI9wI4Qgc1W5ME8620AFaRQLkVYlJcT9BBQB9Dn3EfDnQOsB2MoLw
Wx0G9WnsqRJ0x55d+m/hCfisb2dM6yXOK5SAwof22yp8EH/Ax7v5nQTnHZa0GVq6spYa6ik7OgiN
7DkBsBDcO33UD8a/svxewtb9n7Wfg2yxvBzdFbu/gzbOX2DuIT5TzC/xlgzKGuKVWOXHZotg9k1j
GMmRfgNjLeHeO2z4HgqBPbtLzAQD28fsH1/SsMnH7ouCVDGdGMzSau1Fj89g4EcoPggJVYiRayrN
yHVxFiLcl6oJB+supgnWINyx3m62umbQVlrzOXi7u1ntIz2Ao2vHh/V52DV/UKX7R9rRMfeQy0q1
gp7wKkxFBJIz5B5CuUtDB34yhYJ1u82OV1HdtALdKMMk+yqH4BzQdlSIYHBdij4t74TmrQB+3A+Z
Q5ObHfCIj7kU5WkfAVcSbEPHYx/LY77W3iJJV1R4W6EAuqyG1q1l6nJyYJYnaSdInltyoe4zRAdu
lRW3uJLD1mpJV0hepewDyEvmVYeN17tnFTDiP7IsnFdwWnyzmtOMWIhyu1bqGMQmJnsfaRc/fLH7
8fwAeD/WnskL/w1/5QiMiRrANJalGM1rYEtXSmGL3x//SxnDkDuqaypAqTVrF4CEQW1gFE/uqzVK
wiOPW8DaBCZTmV1PkOM4AQROJ5c3eA8KlMs8eDdEt5pJBpb7FpOktHzfIMEcZNovoP/nYauX0IT+
AtcEnI1hBTHaikIDSYAq/7jPhng6k4MOkYOCazmTWeXydQMglBWqpaCIQXF+0C2bcyyDh2LG7WKP
S20b40p+MaqVLqB2HsZVfLy0UeeLAdCeva25W522mXo+WIdryJLwqo6LBeHaTbR+OCcXM7zsSjzq
j0CoGI28G1KRACdqiriE6wEew2neXYdBPQc08GlV30woE/VTqWdsN/DbLS14jaaEyoE4ncMbdWu1
kYrRI68mEGzL/pVVf9kgZmsn1K19xR/tghX3HQOToxnptDO1Eo4K5DzVmWUCn/lWKE+d9276pp8Y
LvSCw9x/4IF9QvFF0mvGtuKi/uxey3t7evFQ07Qwsv/XI4L87l4g/SM01A6p/huBbB/7D4zPU64Z
Btw8ugKj+XYHqdqBVmuB4TNJxBiJmujWGDbI4yiiEbrI9PJRwl07TDfdxKI0vWEdAMDyZH/4onOk
M3376X7zULNf1K3J5VHWU7z+zKdme9u2sGxpVBR4U3HMmHqCwjBL08hPvF+mi4Sg6iBN3jHZ40eQ
fFUtCpqywc0VwRUiU8/FA8Gw9SdYRwuaa5bNTnKJvs2sNtwMX0iOjzHbCGrGh1nG04HXNhTkeXkA
S9sXslKKIkL3EzYajkfYMjXdKu7IXXfaPirE8dJo0ndqPjtFNZHNQYXP5qh7KxTE7Ytgd5rab+i1
hiEaZD0EEx8Zyr6ThBegSnBGoChDzkEPGyRkUveTnAGJt+dTpVe6H5cI0IUl0fIL1XwJwdLPDA47
cQa0+XQQFZwh6Ur951oHcmig/UA+SXi980791E3b1e/uesHQW80VexSsS1J2y195GOonjqJyPRPq
1+jW6kKT1atdmVJLQz2GHHWPgt9QLFKWQu+J3GHvF0+AyAIKk0bmbyNvbctcS4a4ITXC2LpHJ9EQ
bhv7wEYVOEOlywXkbe+fGo3kfjFwIc7WejDt8zojujth8UGkltPacAv/s0ZN7DxbnxDuDILRQfsc
wZjbHPfjnvuTPMRwP7+KkathsRz+1YMcoBvR7uB3LF/P22ZRwt0+eU6GKUCSJqs5MbNF6h64zXtf
eEWBPdekg/qJ5eU9QF5EpMgVH28aFDheWRCi22y4ewP4hS74CzWXjkxDCUoAqYyAJg2BHBeHEAj1
UvmbzDACxdRahK5tELxvQNxwfqVsEOrpXRx2xRrOfvO2EtOm+ic8hqefM2YEMrxAnkiBYMKZ/AVi
6F+2pMMLsl3rSKlbE0BrpVf9YRtXhy8w69IwSyqr0ZQGQn6aSjUWWM/TsJbiKtAlBOiqmZ6qaSLW
JiNR11uk2WfZluo3vAt5pketz1Ls5sHCOLL4wEdi6lpyG7PeU9OH+7SgEAkgMqfvvsjqzZ7UAfUW
OQY3b08c2ZVKmkcj0xDz8YRRxEARNo+3GMt/+qt3HTcAAaH2r2Gu1nKyRU0mtXMoaCMxuRTPajnV
IL5r19LxUmsvIAo25eyINtbNf3tLzgzFKbcZubJa0HScSolJx0e6HDF47U5l/CQg6RB4yOn2sfBq
Ckad9k0g/wzuMRUDBZpo8zkFnGppOrqFt1RClUQdcXr24yn/N2/9IM+uih2ByFL/SirCeNYOLWFs
hWxDZedH3CIPPLKaOI+SkKqFXP/TDDLyhYC30Arj8DHOhfZY5lpr938BlAS5GXxVDLVxgb85nwZQ
Zx/Yx4CuGRKC99yPWXRRmwdxw/nlFR2Eb4IcJ63wGI4omoQulBgAmJMLYcMYJ6wKWiNunW1BW6PD
H2R/U1H7gN6BKlXwwN8p9gjgkfjfJann0Bt5JLO0vtm32eprss0/ZU6WIS+/JhIilJpBVzUUMDXp
iBN8I1tSxgx/O5zuawD5X/VuB4BqxNSlgSHCyttbNdIkPWBORCfR4NsBFjknwzGvlV8nYonZXavB
MDFFsVsBWWohOGdNi/ltG17kOZZX8Hq7HJeIj0lCIKBjW1/TXicL5AHvVK4ySpePI5FwM0rpuim2
6u/UXlzbmAFKGjCRmR9iLVXWsVQ3Cw/xK/qvlOumKUCRD/cUjrrcYSE5H9P+iad9PTdFH7fvTjEI
IxRTSO+Glh3rt7HulhsgF9BbqSqTEwxHrJ+FgvRFvSKAyvIvUc85Pq570crsfGC4jGT78lI5L0pn
/pqQbOrPXFHMCU13FZl6utZXa3NWhediWY0PxdZwcpXa+JcUtw0vjG2PPe0WqziA3n1yI99ZAtzo
+gf20xcOdSax+KdLFDF1LTE7nrafU9X6v5SM/qCy+uCXZM0QlUb51PqaDpq2Bq9F+d8CmBV+srhK
jq8ZS4v/rL9daxADmtV+IWBvf9NVjEPvXYlAIIs6meVQq0VTVm77ZCWeb0gKXxs01CplM0G2B+q9
NWPQcDuFQQikmaS7ceyJsj/FY/qrN1R8Uxqu8dJ3HJSeqBbAqSrjsh8B90paHswUZv9EgX9h7bVX
AeSCZQiNmtA0It2cDw8SypviPo35w+6aj4Y0D4INWR5dPDGCFi1FQyYs6nYA2o8d4hE8Jle31KmR
cxeb+mt/vFHk/omAN3STfjixsZSQDEJF7NeoCwzRxS9z2Fh6lHyocYNPtDy9OiYaCubkqDA0TqkL
L4ge9XrGYV57S+BtfMcIE7AnDwYCjTSEykrvfcLHOrcgaulo8BWAr/NIef/MXCsNFGHhT3/remXQ
MGsPFQcWX8s0oLvUWJYj15M00wA4OzpMEgK7D246tVs6Gpw8tZxjaLQFntbvtr98D4SDjKL39BY/
PlA+BAa2P7RPs2kmP+DTRmjJaqv5qHsbhcBeB6t3Pvq89b+eimk6OD66aqWZf5nM84FtHpxL+NTM
Iiy8tBXXUtpPCRy8hthEdW9hmO92YUPmwQ9/xvt7QydO/1usNlCQNuufC4h6iIZ2QlONckjojsBb
oWHOtcioshuBDMPCDVLYrODzxxcLIYj5t4FUFnVrgfCh/lOOtR0mBbTPHYWEujqCDoLtD4y1WSG3
JUp8zRHu/SxY1eBmtCRpuQwDpdmp6iwWRL9iEckEQPYkTytXlgiaGEPF+vUf1VTnUORMAleaIV7d
CI9Za/bR8Sobzt9IqmZ5LgBaDg6C+M65RXc3TgqpUDtK1XgtzQrwnazPZqlyPNunMNqrk3OPsbx2
lygBeSQm9rU6fOFc4HI6e6j2tY9iEP8WOc+C2viQVVKQ2wkjgqrOurtIIT7Q6146M3/1SVSAWsu9
V7G4yAbwKcf2rJlV0tghVgY6qWQ58qS57wNVwH/T8sfGEVgbE6N2DCHwr+zy2heKnTwL5MmoGheX
hjZJbzR8G3ry8xVv1+/bGbadWfvQ+N3a75z+1QcJLbB1GhlBJKhoLosEscT/CW/6QOEN3t+Py99c
juozKlI8+HI0uUlxHlW5FtjVRNXqIIwXmzudcrxm487JBoy8keByzt7X9beqn85qStlXstpvcZUP
9iLiAfZZ23E7I0toKlzO3Dhsn2FjAV2rTMB2xVFS5VcbFewbSEb6WpvLnxib7+6AqRCo2FQELhee
aW3v40MACeomHqBexH938mzhrhQe8wqZMkspW/7mO17vjANyTWS9ekkTcPwv0Pp4EkK2KpNI6zHD
XYyORDgK/Sn9oFeSz3W6czTRYVo5+4VIkrOmR7nhuBUcZTkGeXmkBwZl60IGEh2/6IrEz/XdExmW
XaHDlSmsKj+RGWPJQshjm9lLpTeRw/twbzRKkwWIBaAeGUomCb9KXQm3CWWi2lQl/SK0S9Yx6rZi
uFaljeKnmbqJhJYByB4k4kYsVPk88G9uVMzxAVJp0EcgejTa9AaBRo6URqPe2ZoD/d64756NxRsd
+vw/c8LW66oo0V3eicCObzFm11sNemcaEL56MxoPlAERjXffJNWSRCPd52LB0ncJUtVTe8Gt3zLL
FLQllzNqckJKQIyJY/Midp9wVx1s+E5GVSYu+MVbZDJ3jBBOOhuv3CuIEjqdQyBCgLBoKqO6m8dM
9quAAyqVRLYfS2RFDQeqow9hKEWUAgl7uwG2JDNpWTNJ/ABHDNNTzM4ofiiPzcosx4nVPvPwCeyY
0GLDC3dzXpTgKJ5sEzcMc5WKHv7jqbjBoO5yVEb9hK2Hip22gHR+6ESREsnVJA6VafKpOpdZcmnr
sOUF9zno4dUoSVB9mvtCmqhtOMRbcz194yIJOU/7negMv6pqA1pHaX5hS8PrCiouh1xTomiX+CxV
c1h11/FxbDoV0uFtsJWxVCG12YlpB4NLnSVw89k5mo654Ja5fJSDj5SieaYeoh+aHFPhsF4XnUMk
gCMVqauwPKj+O7YRkLPlOoWcEfRYwBKPgzFgODv3AJ51ejI/34LPkZIQ3/dMs7KUH2/D1biwfLEW
SoO1lBW9fxaz6MgjqyY4LYY9FwA1Il3/xVJ0+oBMq3Z0cjZSDmsVd3bHenHOUr1idB/Chg84KDwp
V6uLJrSliWktDYM2vkgUhOrZIcmV3XpEtX/6TGXb6/REyIwRJhjVRUubcYm79uFbWQgqgLFVP0a/
x5sbTSoaSLCbnwM4hGLJeK9uF9XyjgZasBQo7x5i6EzyuAimcwEf+7HqLZqQdZYRym5Qx4qGica+
1VuK3Wg0TzjYnGsDSXNWmLfCQe6tjBY5noKPHiLUNigwhwVKwfnP4MrZRlnMmeXFKZ5/nJ7axory
8iBPfVdhc2lck86dtVtSI/SJgJyPT6qdp52DUs6ZrR/mGaDX2Q3HJxPXd1aU97pEnpN2R5zg6veA
Y1TY9V+kZNxiusg1dGB6Nj68hlA0qoarUzGGtADMP14Eehz+jENvw6clzLexYoQyv4lLRn8kup7u
JS60yUkDECmQGYO6Hbyoq+u4tK/RCiCn7QV+prmwkke5RXAPtah63vsi86BhwtujgtsVtJmW23sT
PxAhXwzkzyL3XohLyZo1SfDkPOaDDggLeY8qbrSIS///5JjfbZ75mSv3ATdNImqJecbfcRRO9n3B
8RkDCih2ih/HPqqyXDCmeflPUFAz2Ngjzvl8Qmciu4oIKcJWj7jBQeY4NxTmbZTFiMoqmR0WVEKN
e0t4FLL+1LnB+v05ul8Fk3vDcXRtvYLAEtrSG4h+yaUrzgc7Y4gOX4fpM770bqUheM1ecjENuEmL
/buwd8CV2ELFdQcc0sjtecVzT9Ic1nS8Rtl86G4XfZsWxHCyToEM3XoLu9fGHmKWStN5G+4deJIS
DZpthjsXCOJwuW3gm3WVlpIvw9uJDfiVOTJpqEuX8GO7CVBMDQrrOjmbK3xnOdxIpgzYCRTbs4Vz
gDhdiPoHgCXF41k7m5PRhUyON5k6lyruzX+6uofY6QTgj+wi6DALlfqqq/XGFzNnsBcZeF3XWlZs
5j2E6YA5epMCBwYcUDrOyTEnWUjEWDIaAsdSHAuyPaxlMHqc+xtNmKeDiWqlxNVv/CISDmrMPlLe
SpKrdJQhNaL8V0Dp7BKVoBTfI/biVvrfh97WMjpKc2IlTOPZsArvdf3+yLjzu5WxEDydSqCVxin0
Kc2UX0vmQ35V91bzMJzB8AvjmyNvKXVy9zSI5gFe6Hv/dOHnwPmhI6JzcPxIWCfC9QpR6fh7UuUu
2OocVzbbaQRKG1N/zXLqgtHUK6ODYpfKm66bGw2Gh5y8ItJhhZTQSgnK1SQZh8ciJ3Dgck/R1tsr
r2OujFgMq3YigZZNj8TmGWiiFui4/Ae3xQ5t7pad/sGpmOPjCNVmiPWMDKQxNTc7GrOS9dh87jgw
uAJYnUZK6D1RvAJb/3DsF0Skb5C73OvbDEjMNnNqVJbJwd14sl9Mx571IHprSmh/c8U7dEPDsGBO
3I03mUNBkUhYX6h4dz0FwujGtlWI1vo4LUIIg1NB1jBtsddhG7vJegBrKIdM0xwG7Jnk/LN4XLnN
6vvV3lAuV7w0vZMUkGfSZ0Y1WaJhNGhXlLMLkeHPqQ/auEtfDeIEYbHMFWIZ/vGL0qSMqxzqPQw0
wCcsJamRZpE6010UrajiMUhpejQojbu7Ccs7ukg59a+uPJr731M0stP/aKL87rsB4/J99K4cNGku
DSS+VdMnC394skCbsuMPYuAFgYAK6D0ChG224SWw1pOpHFQ90ZBNWnu5iIWpc/6UM/jM7ewKlea6
m3ZjIUXcsyiUOD6WfKjpVgu47AfDqy+a1a1/utd2YhL/PM9aXx9PwSRj1jUofilDPjf78nVooiQK
B7MQwarRi6KxOfQXuetMz3wSAthsMgYZjQg7u4HmJ4cnXXK1oYcxu3GgH8W0xro7ghLdaGlnIRJl
f8fRuaYa01r/1py380xVi2PF0Q/udv3nU7DhnljTsem/kyna1sRwz9kmMOr748rjDv50Xavvagqd
xGTf6fiJkG09jkUU/E9zdfkZ2AcoRXEVHQZS32zdQLkLWGvDIlQSb/Li2fMVpApiArP29G25pv3U
RGawS/m5Q3s57plQtQk4yLC2Yf2Pn9KDsd+WrV9oGxxm9wQUFyjJrlylRX/BdG9uR+wjFSHee8+Y
mgYqBAV0EoezOVlSovY3RnSpx6sAzECmuwzXjdocnwLc89po/zLd31sKTzTgwv4FvZbXuM0COcGH
Ly6YjlSOWEKGodAwieFy2UXuJf8pYGCqZV9+XJ/mtjkck98d/1JbceECww9KCeXADOzedJukZ+Tw
1X5bLlDcIABkATVyPVFHqcClt/krZIGD4tH6znec1DowBteQ2TARFITLRAKjAK6LYNrzErBwGiD6
UZDkpnPpToyGfCbSFbkHr2rMH1ehPvTai9hf+T/kf99mjIINEGOnJ4rzFF8ngEjAsu2rJWNeI22l
AXq4HpNBCKmAO+HLseWXCUIzjIRigFIvDJ7+Aujr36bww2Jmw4KNHBuHfRunYFokpi89zpQUKsy7
wULtPBVxQ4ZTlbU0JHLXVYaNXBz6G8q58xFATlQMW9mdLs4LtxHjUYn+XJIY31zQdxm4ILOmVDFp
D2OYJZy2dGcwu97ivA/oaO/Jbh4V7J3KmY+QQk9+UKNI+BJ3TGaLaJ0SHVJvT8rxKEXFJbuBwuWo
EZeRclZugUp11NEtCjcf1J4JkeUQKHWO3gr3O1THrG+SYVaro9/JbBWBYlTNkITqxSzQuhdT646v
fo8SiFzaAAi2cuG0C9GoV7qQaABIRpJkAUUTHfBtsKrcIfsSJ+aEv1DfRSvM0EfLfbwHaAPvmnMr
ziXzx/MRZLpdaocR+niAzbJDjd2QvBjCC5Z/vsiGd+z/v2LPvDbzE54ZfcIK3w/n/Nup2UPaC+xT
asbwhVjzvZB2899klLoegbGlS82GKUW2zDML744tcHukTZIhxSY9YB+JA4i/6xSnXD3zkOeRloIB
NowZDfoolpP7N4F1WDmBCUqW4ToxTN6DHbTfDz7Z/lX58SYZiZMXGJwf4Uq2dc9lP7ELQxn4k2Dt
7YdMle+DYKZ8PhQjUUGWv3vdXO9ciJ2oRPrEpj3pDgG0ag8J1HqGktTbfC5OrG9dMvDHaGRA8ReT
9e7PwfXX4fm1GrvT/Ia3ILWkZC+aPJPzwMrgXiCchMvJs0AbudsuBU6DDHxVwRoXmGQlByLapNIU
XLNHxKvGcjD9oi9ThENStz+OMCDXZqIJtWOVgFhNm3zOXiSiOk74N6FpsmjWv959mrY7VpdlrnKG
b5TUiVCLtn2m+zy3NOOMzgEGo0sROtaQ7Tyau7ZdKBLDjlIyUbAGS29s0q892aZz/g21ToLjPwli
qVtFJIjr7ycDKT1WPxGnS96Up+4BIIzjTZHS+ClbCR5o5kVMHQM9StSpC5+oyCOI0o1TeEWgFgqe
gGYoZewVuPrxeAZxP9OSCPWqPQXfEL5Els6sgF5dB2+DUNWuOvzlsvKlECq1mOZ0UdEXNZ5je4ZS
fWq1Y2jvSsefIZCIUGEmMok5QOiH2WRiV4SE8mkkLsn8eqyZ+Owba4gSFf3acG+JZ3TDPCQn03VF
Khy2Lb6oeH5VtsGkWpvNOlTEXfr9MahSdbLYfM/2Bpy8uLUQkU/sRUsdGfmx44rbG2Ah2d5IqaEB
zSdFGrYgJePCkgVU/upQ9YtdbeP0y96+lISarhkMsz1mrGFDv90KG3eEADqSvuGm3P+hqGoPuRHQ
Bm5stPHO6gvxRMjonwAScBndcMtvpVjwilZ0CFBtT5N3vZ+CQ1/0/H2ZuAJEiOkVwY7RknEwzleA
Gm82LN0C2bKC++Ama7SpN82CIn4/pWLpN08tBal15c3AWJmYHsFuAR2s82RnK0c+bZEqVVYXRS4n
UfkBO0qctgBNYYUWdZeq0VpRtSCrBfGm7j9U+OvRymOfQgEF6xorSTR7kkUCOAsflhgWuwgtpCQQ
4aU9Gg6TWP7GiyKF+FOd2r2KBYr27tX7aXb9k09LIDGngkXlb3KcdUNW4LjOteZoubhUAC1aMZQy
1Y1fHJsj4zsFzVDUIHmC2IEKZ21z+ea23zAQ/8Pp3jOnSzFy+Qrui4tJvQBVCPwPYvoXGK/4kUiq
HyiAsv4kBX8wnrWTLkRNYtTnLRGNfN+lx0A+9KkZxde0r9U9L3ZmX10+0B4pHT1adq+vsCy77/Hx
bIMDwaU2egWqhPm+2ZBjfNxCLhsL8Duch9CqhRg5fAtBmPgv27+Xt06jxXHh2oLpqCIl8rje5rq+
+6Fi4qjpxYLc8mj049gSVMGsHLn1WVv+hLSLlXvcTY0YrkxxVjCnzgvCi+q2XunMa+eK9OnQbrX2
ExheNvtmYtGCLCLcCd3s+thdrGSoUnTLkqkWzoz4EICItTYh3Ll5TliA8HvKOXcduAWEM6U+EEnq
eLBTXpLSAtnTLDcHsQA1pLM2zSNTwDRqG9NcVXh1RtR8HgxuYvyJnvvjtQk6ColREsoPu6lOFiXh
OnipOn9T2WOC10FSP6Mj0EmWXr47QxjTvc0MYJAayz1WzVUPmahSPa5eOE6Kq8p0TNSKZHF2VxKe
PiH5MSluXEFx5ODUE3LLObeJ3xYQkMSv7AmssD9qcshKrvBLhaa7e0KoZI4zNSzYgdj+v7bgkTKV
JNYfK1epmO1bTuRv5Bs8lQYcXWYWtXtuuo09Kes7csh7pIh8JZBTYjF1URD/CY40dyTZJemNZxgO
ONa+terzdGEVVpTJ1ajfbXpOzH8UkOWGvSDk4JbfhR8BfL5HZLg55CmJ5Wg51cb1Nyhx9//qb63W
ZtBDxZNEHPPvOAQgJZHuII7UjXmkS3j17ogBHqUbS2FZKH/Noz5UdB87FWQCzQjkNJ3m3t0QizmQ
qhXCOdqO8kBadYwWGuEUDvQ2yKi/8MYrQUibOF+7i/x/NvkYVACo3EP3naxC0sEbsKeSVWokf34c
hJSCXw0Tg0HR1ritvIY+W038S6n+oD8EwJMWR0cFrYa/fe+N80O2lJq0xqReqfzc5RrJ3s9moK5H
7zVhCiBSnVNsMSg/DjhYaZlyOEidKAJwhgdyPo+2bgXaq8Waatrw9vOFUQBRy2haMcbjmhsXiH3l
epPxiDpPYqiicq/jS5QhtXOmoOvrA/bNl7kl/y4DRSirFA2kx23LV53Qnxp0+GX1dQY/AaDlsJe5
d5Wje/hMH5cJ0rPcSWMav7WanaYPsprz+yOQE+WzsNyIHDV14Z9L8+IaLb2I9bfRmVp/wl38ExnK
jmM3gRaeZg11WxdJo/fUxArOkb8CC+0a086oXpQUKgZHfkUqzUToVCylp4N3ZuTrCxkT+V0iR8AU
fzfqKHAW0boQP1Gd4vs/UaWKO9yojH08FWJCoAOWKKWqBJvIfCCMCy+Ldw0Z2L2dRDRl8sdpHQvt
rC8DQPp9OqMkTW2f7+xeP4N+zLx1R0CKrG2ldSudizb2I7UbD1DZnOk3AbsXyWGzFzDskbRGCZnF
7itAprKDBhAstlWwBdtfrAqCzqnuR8xQEvY71SRFq2weWUOO3vPm+arAB8CNypkPpBrAf/WUXjMw
5q074JAIEI5VLTLIydmKrot0/5VP/O0S/vnePhxr/vmuIJ6jMj5zzBMV/hsvoIr1YT7r1j0rgg4K
ct1JjuLJFLGmDzsdVM2M4MqdHxGzhrQFgCU3kzTkvS/pvpvJ7gzS65IG5wdFRuqa78nvl8vtCDrt
/pbRwqbwlJyT9sX7PQKZRcYd+2Ba7lQ37UlvE7bwX06zhDPtqH58b8pRILx+LdKBLTwzAEuM4FwJ
0HgVdVFXD+f1Y7p2dH6vY9wGqcV4bVVp9iODHuYmORPksI/kp2MkJDcquqLNUqk3kiLY02TSYOvX
EAz1Ez3gPJeBd1a4R85lUD4+C/SWdglNNgV5RLD2ob8ZCQnCgNDLtgVlRLXDY/JyCSNvHrf26PJ1
4c43Z2hY0txIkY4clmewfpHKMZwLl/YVoxyiM/pJfN/+y3Gs/YkWt3cIjaoyT71xFtRLuezI3CO5
7lb0EPs+qQEswtHHg2DYgDoGR+zxLPJOAjZR5LmZcNyyZrcwOaAN3fNHNrv0eDH/KC5u1KO9hM3P
BPfv2P7+c+cr/Y+2SL6wrT2rocmN9BK2NWDyZsdGwVOksfho4VYCIkUGABuRrbpVoffM1UV8ovD2
9XM/0KYeiao2U/aQFPyvR5AdKehpMet8Ofpg4e3aKJdBzFlBsWAhUr6MEvJvc6cyodoItn+xtL17
gRWNLCX7v446mAVIEld9oqmKi9DTuzhStEQFnu221IJOTG5HlqTtH0MtCMMDMBNX2AL8fET5cwVU
9U8IyRUcjt4IZHY2Vjah3QmlxeelomFvkFJHlCQDzfpJbHE7A6Oaye/x1no1EB9XLXktohneTZrq
Gze+iu27PDvUr1uIkJQoPaT+enPaRj6cQs+/TURMHrzc6WA75Zm2y8pUAJcz87q2cuDslgCTOxDl
5tzYWs90Er2OvBLVBtretbqoyN10sM/DwKr4tiP3PfH0MAcOtJKikl2jdU6BRp5w/Rv0/r3FSZhd
b4zdWUpCDYQBSsdIG/qIlRdE0IpIhTatO1ga5NxoyM28m8CwQB2rnNdQrmh4uoRLR34yhsISv4ml
zxy6AXVcF++Lwj1g/SjuqQcuZg/ZiL5GrPn6ThTWGQ15ZGqJfJHMTliE3wBYUSuTc5Cb+rS+u/ex
aEbt4R7prrg25mFvaC46NtTrGl8QYBGcXVJ9zoBZWaRd60yEH56iyh0jPWsInu27oo0OlzFxKmqw
s7cPKJY2TEcOWfaWoF/Eb6rkXKRCPy8terNKlstmJ+wyWGEvgYjK0EgOAugl7d5c+Mc2cDAkwOlR
lENMuYq+U8GAiTZGrBr3mxpW4QU9TSJnc+D/iX5XcKKcaphSG5X78x1XNKX9tXMvayXsGKSIxSdb
0X0088JHKEeRekvLXzG9h1FeLANn1XdjW1CMhEtPv73fQovvqQkCmITWOROhOdIKUtHGn8E8eoXo
o/dlHYLG22s6b7wOiljzh+tzksxb2jGJii2dL6iOhvHoe2pad3NxOJSBJ4yWBiGB7qT6SzNBB4oK
FraBxqL8UduScc29hObO4U94zzt7LbOK4RW+BUJP2kVifG9LqaCU0QnFKmu8lOSes5v4usVny3Fg
mbNUSKY4eo8jOCaqrMdgl6T9qS4Jqvtg8Cg6ql9hMtJoi8I6OCA7FV9iun8cUzPjMYzmqNDHAMpX
YfCS/j+s8okbPg9HNlXj0K2ZFGgW/oojEVi95IO0vw2NuTdV7lTI324akI7VWGjws3xO6DBSX54g
XQ6Bn11l+KeC23q46WO6jY8/ZgS/F2Hc+s7kGAR7uDpqJ7fzRJKQZzZi1gKGunal8W1f3cm8DBmo
qL6F9H3oxqnGoqwgXTpI0GiDLyWjaQHJU3LabaQYQ95tyrBmmAYkqXh4xkT936iWPiJe3pNei6LT
/80MkAx1aXHoabVtPvZXdvyVHVx49n8d1WzPcU6iqvsx/qre/bTq+dq7Yhn9qLWeC8YLdhExXVQ7
0F5DXNTBIRKavCxgKoop2px90WgL4PNk45LxM50R0hmYd9L4N2L57EjKOeuPykEsZ6Eo3Aonvf+9
yOB4SlgvQf6SD7fS8P4H+gApA+LSj+YbkMUhNgCW3rZDU/rV4XpS4hIcBCPRshQoxRim42tLLA2y
2boKC85r8RWvRex2EGCwmUxu++QWWM568aXWqLFuJBT0AycFXQJiIiRpCtUu1fU0mst4EkxIn5z1
1V53ak3pnQq6AGwL5YRBBT/riuueXt4L9EOM5XlbPCOzDZgYw1VOWIdePagc6NNsITEI0INSiX0b
ORD4+xLgCrwbaZQM0t3GT80sCMdZacZdk7Z9WHtfaQ7AUmbTcK3tFufDhBKGG48IIrdTZ0ZGjaeA
4sU9gDNTw4LhGVjw26V5SDvFLKFmWQpzp71AU73sfWgS4wA/e11bNT8crpBAXizf1/Otzkj/m94X
1Y7tdjZNtGmUxSpdLe3dJ5dXOq/jr51oJktbjpMnForSQB9N5Y7DTkGEMEKH8AHShVIjVW4Qe1yY
ZdQ0KowAJU7/OB+H4YXtcGoXGLbYrggwOpE14xyXqeB7y0exa3m8QtH2yzfXM2kOF284SpDDgrvM
ei5kWnyMpSLrtsIVoXyb7VHE6qa9kHGT6jvfNuhhlJ80dcg/HIZx7M81KOPwpMN6t0oySozykrO7
CFbssZ/SRSAD0CqQafFKUabZ02YdvDyBh567GNyYwtnxVWN1/kdpuwwx59qTXqQhtdE6A6PYd8Gi
4a/WsE5igg+sBvsap7mhgQDmlHss3CaEW3oBciD2C2H+sWWT8MuCk7MPHtyGr+PchzlAweSjOoOP
AxCdgXY1Q69+hOnJS6hStT/qny7CCaOQrZVkxGMDXWV+QjIwTH985forUSN6pEdw0HujIlyyQacV
SSRs8O6OxuSgqY1zHiuzAKKR9dXrV06ce6OpDdS0yzEwSquyn1B4VfcudZIzTTlF+ulDiS74iTRP
XaN1hTmMseb59Hlp+mkv+4/M53uncZj0HHlUS6zC1eujTULueHxp9BSOP+Z5BsL4kvIJOgvqWegi
XxfysYfRNm66Wx+WgtJOryMbUrPYwSs0nUQIg9iS6Fsx3zm98gAL3ASCYxHD35P4EfL/0FHKC6kq
N8xX7T74DYmcfzpaQawJUyaAmMAIuOUqWrmGSy/sugKNthiInQQ6S0W/a0Ncn76N/ZP93PGRjX1C
++5H3Q36vFsfcssQ2kFO3m1en4fXWg/1jVFHdoGOr3DWxz4ZPL7guRxdmy2n84q9rlqOepfVpX9t
XEf5xNLufb8O4vmzBjMtYC+4tWzHaBma2Es81m613ThPmjBjfyS9++lFDwPPGTCOYC1XnP5Ye8jK
ypYti3e87SV17geuVD3ZO+THccUQwEX5rddTu2V+Np7IGXyYxTLpLJzXQBDskqlZJqd3nXxcEaP6
d4nE3gJeu7IIuP4DJO1yHsh5oCRikEnYklUt34Lua8ezluPv0OLVIbSiBe4k29ez8NDKB3ta7z7K
MZSBQpXsC2fxf0NfQwBfEkF2IAZfoBCOaJJ5rYbPhZaDDYxYpoOOHV8JZNlzQfg6MOi1e2r5ZxIx
JFCFg/9BgRwIfjCN75ydz+E+FRCgb28mCDUaghmLcPJ21741YNpu4bBM+knb+fhOzvZRotKBLOBy
quzcG7lMsEARUqWL/hPBJ9Ldfh1nXWf8rEuXWO7BvMANpvHwglgkPI7HjS9w0ujk4ZVg8vw8tGBe
MYKicakFkYCE3YfXHklPuBJIE5GfVN5e8lflcAKhIieTj2JjdmleNnAxDNfOB5dK8rBF41V/n6ie
47q+Da5Tl2XvDanGr/QLq9EQhC0vn+P/IS12bZdIZCSOeT6sEkrH49qLocaclEo/8lxq4pbWJ+LF
JDf/9ihz8/wfpp/q+0XqYsxXo4D+7r+BnELPoXeA/VxEdVAu0YXmZNt5/WjoXQBlv2oqfux/Oo0X
LysF382PT9YxbjxadW/k9DUi58RGjunu3caGa0ktY/pThI6b+NB1YTiN6aEk2ynt7m0iIJpDIzPD
uOA+Po0ROeTcxthgkZmSwa+6CFlHgM40LJwuffEl+9iEcTltoLgwdNINHk2zHfnpGqEI/nnWYHyn
n+CWFZZBKjWfK2pMFkzSDanpsMUgCHuFrCqn0i11xelocbh982dSoqoVe/BDUv1SEAz0F1y+rdiZ
M9RBPRlnPw3vJkidgSvGHHcpE1AY4m715RiUr39IR9NmgfJv6A428tPieK75sj23S6qyi4c9mzba
vBzA7NlYct/DPAMCNoKRj5lhXVxxMDxlhO9USZ1CemG4Sb5TEDA4MqAOEXJjEoQOiTPnJL8nYI0B
VvC5hZUKX3E1NE95rIQBMGZGhYtpuQeA6iv/PqeBX0ckkY4RsAOimhnjmboAK7EBO5MrxoVQI3Gg
2B470L8uSI39c7h48u1v30IHTSUyqt8qqnJOcwevuG7Lk1NvFwvFvXDf53X9v6bx4/RwuLv0om32
44JaDAyV1Sapy77AovH5NiAeeKMIWC/rfW9hP7qDTC7ZWaw2w8OxuIVhsE4hU80XofMxhqMWWdbz
nxOf2qrkazOzDSrLGGk9ODIJ7qUmUXEwUsiK2SviiRbawlPsf9Im/yOMr7d5kQe5hpbmWyD0yDXM
1vOH3gtTPblj0c4r3uuyjNXDnu7EMcLbCKVyvZhuzzATprULRpLNqdfEGCFTn2bEQecTGmeQcFMI
VHj9Bc0cCKbiGdX8/2Zm/xzsMw/IWySa5VIAzf5BwXiJEQ8Bgj9cfbU18YE5hM/thOpKTA1Bq5F9
vXn2vuFx9bTfVSIar6sQTVMLliUCRtH7CNnYaq4+dTYus7+SH8mxa0XXvNdHT6FQQRSqHRRst9W0
Ix50X6kxs9nbRNNxq9wDktJ3amXdt5zTSINRVOmmsZ1Xe3/4mUU5kgOb/V2RuaunuYW92polryVD
jcteYqbxxYT61mdgQjdY0IEArBnqMqOLcH5XtIn6OiHKDWekIj3x9xs7sJcepZXP08gGHqh2zKMf
z8awOiKVLTyFpESEhp+C8MRZS52KbKJLvyAFzV7iJuMTk/TlE2HkPbiNfP1I+7YCgnI+i8f3qkTC
Es3Oh78rDyzhtz5noXgeVK9gp7CYCUyfJ/JNlek3DfLhWRxzbM82M0+izWMtDI1/Ok+O8Oqbd2pt
bVJmtGR43dadO/iyKWQrIEhxbdSqXFWXScUQhKVWEOc/BQ7JPMN5Q0SDuO+Kjnx6tSov7yuJbPnr
yWJkKDI8vvyeR+v6WDKrxmLbBacmFeQYbGIFeXcvHs921uTXM9gKs/N/UuEw291ichONv7kYcV/l
Cb/U4oWN9ObmnM5uPwJttoVSwivqpGJNSCyALyfyhX1NUzuu+w5675mX7TnSGHPGdx9C31riBNc+
YI+yKVu7fZHnxl4htVRpVmj0X0ym1KwSWC6T/03W6Wl3bLRKLSsAbGzWLNjgD1BypjepDGj2Eh1B
yV8sGIF3PFYxwCW5yFla+3M9VWlUTFIu0tITb3fAnRvt3nu5/BwvlG00BVwyEEPf333wAAYA9jbF
fPi9fz3uLyw6yqqQWQDXsOuLTI+vyWAw6ico0XcuezuruTwRJFwQBt3oQe05LHs4qdA8v9OGMKqP
dxF+uK9NIvzy2GTNF6y11C+GCwG10QcCFFpKGB/Xsx+gFCXPE0z7/RQ39aafANLvN7GPfe1oKIxP
yhlkpizcyLup2mNctf7xzf+IpupwKyDjNNE+uqo4MagMhPC7fX0DtZuZEnKmD7oWNH+Jarl6gykR
nDtzLKRaB/5vLcdBxCEFZoloX2s/s/IvwRbBc9Z+QEkZNJbQSrpw9fjfPU/TBjmYVPN9wr5O6Ke0
kfjCnGaE9jmdUc9iAvq+NzK85N+sBVqm4DAMwhmazMlHxGV/lEFf88y8zALKxSWNEGTCrvdc+OBO
awnP9ityncfKlELzVRymopuz42cxAIm4wDxVckay3rZkFAOCJKbFMjnIakdG3aBJYWCJzPK1r0Tu
95OjSYLXuV9LFxpm72M+7kicQLHqcC9OROASNEZ0bYLgffIwDS9q3zQxIUhQVsb/agxKoWGtYKnw
TEWsPFI9i8UltBeePmld+yRBD8FqTDBk65lR5uOCRPIOeOlHoq+aw7Sc36nE+H7Th4MpzClNhD1R
h+HgrS3+jLtbhOYyz+EazyaVI6oIecBZrCVDJxJI5rP15YOZMv1UV16w7PWXW7+gUdfIxKs4iliI
TrGeTCIHvy8kGerJVG2HiLn+xpjHqhi40Tiqb0BCivmhCLkOUpM/itWiCzyC0E0ycT7ktFExV3Ra
PUPwm9BuUW96YIrawoW3oZli12pet3NR52lH8rqz2uz+p6lmn6GYWr/mUuoorG4ijAR+jPdRT2Jv
tZu+TstZlQePx+g3VUXgoLHfsvF6NekldD3Vgo/ReAuzmm3dgzkNKqmDLxAEMekatxeyy1VAorZ7
ihHn0sSlSPGx2iTYzOtoRfcf4Kgbh+oEStGy+FBXaWqQi7dU1FAV0/dSBz/a11Ukk19JvwmwOwQQ
RIi6f7WIJB6PVW5e0u5uvng9PfQwhisCAONP1zof9S2vCBsQUmb2ajIBXByisjPke7R3OVypyZ1l
txRrD6vmpt0AJWWqT3ZpLRjUSHjcfmube8zdZUm2LxtcCm7HlzEdUqyIR8/M6qZdiRu0jqMRkAWw
xh3d+UUCsIo9XFxOOqlCCxIoxAM96ENghIH3WICqs6iAMMjQCPp/PODhf04D3gUT/0EeUkBhPsMq
w1xKN1lLSmwcpCr1Zr94d5F8adXpsOZh+Em6uGM2x0E0P2iKqvGwKOWKdjCPA18jwX2HcjKIW/sQ
Auz9wqyvSEpL3ppEZd6dxQbDOoDX3W4mkOYGl4uSODJaQ9z6q2YvA2eOxB4X5sDX26EL5JHIe5h0
fTZzCvK69WJgeayJk9A29477RlFzcYIDv2Hj3puAS1H34T2+TO/3/f6tVzaoFricjaFKor9jNI4u
Ulfy+XvB94FDRWF70VmdO4M3g5P8AnzOJU8r7u5UScfqbN2n3CBmzQvVeYPIzICCF9UZ+tj+zY74
OJkIVOOh/LEO09nZ31cGYgxjol1TP7A5FGmZVkmknebNjHJfl1v0VCvylFJ3db9DYpF3zuPdk5Uw
i+1CWhRRlpwAb7g9zWbGf6iCC9EnAH98/4aQgOAY7dJq+JU3AEdQKScoiklRrUHBeOi5Nok0vHtF
GQcu2jMM9QjCnsOMIIRaTNPmVxhNv7Y+Aly5b56S0dJh/idADNBDP+YWGYzDtEdNionpw2hQSjfM
lQVSXu2LmpsFyxdGHOwssTeIVx2GgxxlItvsZ9+gCultUirM1fzAfHCTetBAb9FgAleitn+SeaSF
6LS8zjVO5WJ0SafgF0OCLqtoxG2OxN4hmrdx03YnGW7WCU5MWjkhT9W4kK0HvssI2J0/Zb1zkx41
1BW7UIohj3AnLg7kLoazzMHaYcRAWpOlSQOUEDFH454zP+tTcXlgK8Eu+V4QnlKbqmBu4BQvdhYx
vn6nBFX8tWH77nNyIsZyHIR2Z5YG9gXcjm6Yic17amjqiujjGao0XrOBC5QE6MxzOWnfqRxkaEuh
Oxt8PtxlVo1fxSciL4YrAmHIV3/seDTRgn+4s6RFyyAmBF+CgYoySW83xcO4DfiKavAxOm+/HaY0
SxS88F+BzCCVs+D5Gk0JNht7T6kkdWM5Se3VpXHbQomnOJPUsQOcY4wUVE67fMr2FkLcuDXdk9t1
tCJXmQaHtCctLEq8Vkj5AzSewbhu5szQxTeApa0WzidIqUMdOxTH0ShzPHwapJsC45S3uH8+uSTz
txYeof3MAizQ2b1Sx6rkeaXe6Dc7BwKqnvAF5l7+KO5fJ2BI5RXzr3FcPXh/o6yEdiBsPD5FgQst
7eb/C53YMsMqIN0eoS2uXLBIt3gwmRLTJMAwB5VpROpVcSevn8IKPUN2bhBv++nFGZ6qLp4cDFoK
EzRGr4pUUwEXfZeGRu7XjSW39E6HjrGXYwVuWL5Ljg8Eh7wOWa3Yesl1Snrxr/fzMZr7768z/vFa
6Q6cuqCedwccliHrP5Z7PjHU0iGWqVDNySb0qUAmAeMSEnU3CfN9pv2D9BXTwYnFgxA7f6VJ1mmC
hnDa2OHZoVtN6tjrXb3ExEKVQbWTTLcKHxQ78Vb3BjDj/FHhI5kAH7toZAJ1jNDosovn/DWhdsgL
wA5VdbNmmDaAZnzkH/6wH/pVPphQtfmMWmyPDV+zgxwKomtwWdid780FHOV3a/nm7jKNJq7ZqdnN
ZxOMhZKw2Q7BU0VeXQTI/qbAjlsFiByd0+Ufu/VgLpCYJ/SPzu3qSHFSQWRyRcRx+vac7NKy3GSA
DYxJ6rzPW9JgL4TAwMu+GNOFbEe2Xp5380KpuZXTrz4rCl0jKUlT8oq+wrRKRV4Zk1jxqYzD7ieV
/nOY9IZK6Oi0l1rkbdVsbHIZzGZtMpCW8YFFmHbtz1ialE5cSImQYYj1Rn6Xdsv00NnEFB5Ymz4G
1PywXk5k2yyo/S8Ns+SpZYCmBN7KtUM2LVab98p6oVMc8VsEaNWokGnphqkwB6v+2eedORslHTWP
BxJ172d0bjypVki4qGTVPxoe0XtOgoXOYOWgHllf1rg5jn7ROmtmQ8s8TzUWljNhQ+cYq0Hn1x+B
douPqhDm100F1KLOelr1WM9+R41cEwlgCL7j2CVYrrJGB1dmgAqlsFrsqzmx6ObsJxWBvwj2fKos
UtXzP5iO0Ru96tesmsj4bZpm7APNsMRDIPlb2rDeMDUPF+6xR5apvcWlzOp6tNqaKhFjhXitnYUf
XjPaEq+VbmGDWlfVe4LQNAGE4SqTH1bSSxLiPOZxyZ1ltvFsqosjgNE4obTxvVGvozgyCogvdguT
SYA3YnbgKR2Gwp5h3VCmmwTfaDLnxWe/dTcvErBlsacu1qdYR7+3aAQTWmUaqW1OzxSi+6UTsNeV
YQNH57aQQ2dLUnH+SGAEtNpRbaZ6/8aWl+gymLChEbEB7sC0rZ4JhY+nt+HpstC6fGD+6zVsyFP4
z7oKtjEpcDsETvg7gq7pCkQQYiZ6xFOduvHcYVMezzI36SepRRE40ty33x/dVf7wcwVdw9MBJpA1
ff2ESJnr5ky/glnjrBQD3zetFlfdzxrpb9QLEHjeaB8NK7gq2e/MWVcOgMBlOEXfVxuypT7byTd2
85MewHeGk1aoJF8g1As+UbgyC3CThlFvfGvin+YX+UgmP8JGwBg/yd/iX4ak70Y0omvXBM2y2ePV
BwaHU1z2EqDv9siqa4Av2Ot5wpEPQfclQWBaQ3KPRfE5STMgzJ3MbMVua7yF4KJi45rLv9Ylyed8
kGaz5sUhQ9LO0l/ZaChjFrwUxZJWh59dETuTpG2zN15GODcHn+cJxyKqe37yyfhYJxrNueVUis45
MLjMI0DAKsMCsqSpnpoCg6Xrxp6WlxTV2vlNefzWKq1TsT2vYM1OR3Kyt39P5IzM4JruTGuWk6GU
ICZk9tEbQ+pywT7U/657mY3NaWDQnPuvG4qxViGVJfBwLHPD3OcaZnXPgS1/C3Bc/a6O3yj8d2Da
L2lpYAQXCTr3rgtk1SQT9OP3L7JQbGCNeA4Pcw5WcJnuJpJVuNeZVATW5ajkARBcYyc34MJvpGCq
nvs4RR9BvPMItGiL1D1Sg+akaUuDosE8s4IaECpAEpS4BGhJ04UTQkoIliwu2s3Le5h1guGUeSuZ
vAaJ5dI5TU83urm8/gBp9wj899+khHUymoUIoVb4JlPrBKtmTIPZabIu9Z/Ih+M3CLs734y1b1cp
K6xP6f7dQQZANIbS12xwZEJjRUgMHfae1o6jXH2/n+7AGfJ0Fr/JRadD2AvyIupzxBM19zIuMpiu
X/aNcpYQ9LY0RVMLe2hdyf9DYZNDNG7MEUBSX0oSDYO4u60O4h01DeXL3fu+lRjpkY0sch9mlgTn
RM0YQ9cxS6AD4yZjzsP7uV7XZoRub3rWSXmTGxIS7oYVwdTDvC09nXYMrC1G+wghDFS/+Q4pKF5S
/XJ41hmKHAU2Oo084fIiKPHZr0gmLegJraY+MOCXSIHhoplnzWVDJjiwABvJqbX/Pkbkywfex/l9
E3AgLiFnJxaxibLFpp1xmAjONZUHvK+jgIRJPAsH6e9yAbhauXkhQL8Nf60pUopNVaJRoqbkITQS
u6IRZw38ovv1i6Jv3Slzpb5x8jBxCETisTAUi2hcrBHA8tDmSOmbU72199X/zKso0u+MSyhE1je7
SYCdxVeASHP1pnt6RjPr0KqMRP825dxQzVsbwKox9hsDHhZT2Jd7595+RkNqTKAd9KDiy5ioI6Yi
Atzh26T5YNDnCpFW9RAI4v+4C8+r42DoIieoe9NmSZhbBH7tCAkGxFhPD5NbZUNcFQks9WDquLI3
AZfzhuMyovXldDPNsFrBJqayOZotS8ZYiVHpNDQlnLPxWvV2/hQMjWjfqH5mB8gdXYHUzcAN6jgD
afFgnxk6E1TuAL5HcyF6D3UNbaHiVlogEnB2Xc52ayt/fipsIenwNjve2SwhUjrl/CTNb4NlVUOW
eayyUde9ipmN6F2WXgk2G5BRAUGYx4cDPG/CnxkWZSMfZ1YFwTxu4wGtjJeUpJKP0ehdsHnA1XdX
mA+bUKCDbkgrCe8hjRt0JB632qvh+JoD5HAmaOpFxnGvVO/GUdB5V38i06m6sF+BUeVlIRw2+Tip
X/uLvTIjHSp3U+Q4cgldor5/Tva9m0X+V9p0CYGEvnFSPE8vS5ky24bQ8C6PXUr6eYw97oegOjxT
J/wF7FXHI0fYT9rF/9ZnmY7b5RNhSnxpSiI3t6S2/c8gpERk+UCkdJCbxfrg+cnqBMXIG/w4K6uc
1yh5Br7UZ3GGRklIWOKmp8ChJDdeknz1rZiexgGLUY1Tj4KzEv6XInxY/pKUlC7KdH5PihaDNNoh
ZpstPaJKW04R1adYLNVKODqloGXGdpba9O21iaQrglzowAhDjltVSiMZgoHentiZzRCoDlJi6ygj
1D/M+Bhte8QUfJauZB2zAifKlzBL/fSTkQVhVPlR6aEpdsUIEwMqgrV5k4ytL7EAxbKguEkYQAcK
0O0Rq7Vg0QsFIXJksXANtGc1FxzH1SmFzWUhqNF3W6r0BfV02InIJP/iMWmk5au0wnflgq6Ckwnq
vrAxHHhbcsNSBYLbanRlAd3C9C+iSRJGdcqHI3CWfz2OOcV4bk18hiQKimcLYWpQFyoRHEVpTrg5
DCcAw+cbeUCLVIe1KxJ9C+thCS5oRgQgyB29MaYIcvlt5s6oy9iEF6BHxPpQ5ozamazFiLS7QF/L
Zl/8juYBOQOljqmTCKbvJOal739Z9O4b/qWrGgkskDpvVosxWJl+C6AGmV0AeeNpVxjFHoC5BkEF
YLA0m32Gohld5KAS+KDqHht0HMOQIktixACU/nBFuceXGtytYNZhjXK4Pqvp84a1dIiPlN+RAQ0O
QdsKJFwLXpvaTVbF8Ym7PvCJA40eedwAMTiT+modt5ZKZ1Ge3/QyhbxiN0T7n+zEwsmHlR04tE3a
jtkjFRflBra19mfXgC1Kv/x385Bkyg9fnOQZa082H9XVz4ExxkiQMDcABc5G0XNGpo3y/bTXn3Wu
Z9NHKIJyF29bjpJUt6s7/uhVgk8IqIPNusvIKFtadTnXSHcDJtOstc1QMVAA5Xvr152Dxz2GWSS1
5KvV81Nd76bdMtHU/nc7u3HfBnrvPRtJJsDfYcDKC2LtVzDqIxUkgePEcHxZWftF04E6KKKKCNO3
MELKikLWF5zkUSRMygZNVI8QAm4P2eqZWnt1T5R+PKPfsM08xnXbqXkQ+dJzu92FLjF+PUccay7+
WbQV0E8Ffvfn9cIWWFHVOKBpUTKamvCvTJIkZPNWwyA93MuIENck3aKph+3zjwENgmc+IClL/RZc
GdgciFLfSJqlm7V40jJY2H1MD15jJHVElNRbAUzdq2UuCv2aEUyPls/WK7nGqaGJlaYGq/BRzbjf
Mn/KQnaYNqGjmaK9f+LgE5wBfT2eNXfsaggcTTNngDgLl98rxQ20uV0rNZoP5cwqSSg/Yl8cXRLY
7r30DpIJXpiSMsSD7cjA2k+Xz4atyuCKoYQ0U6+m3kl4w6uglwP1kQQPrgecVlkyaGo6hF+4tM3n
5VBNR37vTkWjA5+hBB4C9G+z3/eQn3h09SXzpgpTVS3VsbDfbQhkDdhH/febAwWVz+sIJGRiMK66
JmbtkBkPjhDV/NmkzekmJwqCNGH4ibuuwcijVaJppuhBUV/Xi6EiwRUDiFiY8tOkllx4ysQr7rPK
uaJNvIXhxrdSu2/vAq7XAxj5Wd92wie05PteBOP6Cl39FIiVBbdZagrNcOqjFOzNi5vcHYrS/7C6
xpODazGZfupfGbHFoyPt8/sycTLnb99xKAcxHOdBMmZRU2/vy8Y05w9sQKs/0e7ALlbifBLpdRiY
S309kD6WgMn/DXyryzx1MF9dOGu1Qvpz9/ezXyF7BkYy5NBPF7dM/BDrCHc4G3JXVCLCzPNt2FNi
CPIq5dNmw7O+L/YyWJ71LW9y0qsHAEjoAs5ugtc0ObElCrXIufpy9IIntJMJZvkWwoMdCRElH/9d
0Ari1s7KuI0vSPmFtYRX3oVy+ZcSSjCenSwiW18fy+nVk7ltHHtDJ2Wa8Hj6Lng6QObxy3MUn1RC
YnGv3yPg40jFRhau5xJ4ZKGis7RBq4wpDxi8fb2/l39bru8F1QjQT7ZFhejWOfGG1fGQRfPHITjl
M2+M0R4rq7Sw+E29ehtmQW8jDWAb8rp7+KMRQJPD+krKiPHRtiWFfM+8IyLc0fwKysNCM92MUiBC
6kA0IMsfgjmsfDHYBcmCDXoagfQ+oob01Qlim4Rj/npcnxukUuyQu3K7TYlxFSLwy6bfYfJnm79J
tY53Hu+R0wT37qLYVJ/M25wL8iUlO9mMSXupl808rCr+B2LhtJPIXuwJ7lA0Fdtw5mwUp/ht6xpM
embhXtE/M+Is0BQLdz7CFo63tuL381dvUK4/N+ACHUilGPACYX0btuAjpTL1tOb4tpuNu+gLyXVq
j4D+YE5jy13jgdW9jXzNhzprWaDFDJL/BxkoailcW/LNv2M7gfxSZtyK/BjGsZJzbZoMBnu/Arp7
GwJNymfuYx+2ZMabpJFRLplyo2JMZaz6yw4w01bzDZlael+8J+TyJN+2xDZW8X19AdP8mrgN3OTm
cpQ0g3Puu/nfA4LD0YahDQShgkrodq12lFaU7jpkbr+sMeoRQTPtACIRq4u/GrbicW/9RzXyiSUz
Fozfmb+j/OfBQZpcZKPKwGYlPnsg5IGISHMQVU7ySakMNw+75Cy+BC/GZeXRLa3R0M9xsQWjYzoi
9IalqVLsYrxmYmY/Wr9hcwUvUfoR5yeYV4N1RudIZMCgMvJJ3Nz5+SPG7gglEhZNpzfIGu5QExzn
8z0XYwnGdlAamk77SkMkG3gKwlIpnNXYUydIdYmeuYnTcX/j0w2YT4/m7+O6SJdIwDPdEY0HNDnR
P7Ib16W+dtTvjEEFWHiqWB2NVB+gifDQnVjAi3o5bGg4AlWW+m+0Rirc743YI9RI3eebqUnctXD7
Z5fCMrI6Zqhayl0wojcog0ssXKmDfOKbs8XekO4sUqGAdqkXkYeKm9ZBWLFwq2oTDlz3vitgVD5s
LHKqrb/4HNbKfCXLHHp//vewpgP+mzSCDN8+k5x7wLcqiOhJJO4QUM37YgxmdUY9/A6suvDmARdQ
s1On/Bn+rg0W2BGGy2GKU2amYNejhBrxE87Jq5B0IHedgdirJgZ6ZzCAL4cK/KXxRILLb3X308e9
8uYYJX7VV74rEURMqfncmcOGjmFhjN/JNvcYKkXzyNVQWg8ev9YgkfYYQQRr+bfo3/9KLj98bqz+
959Esud/+N32suoPH9zU7TtKDPqTvYGUIBcUgiscR6mfySy8sZ0JZPRQfNiUwzXGJQyc4TPwYzaH
qH/zYbvByfXpsicaj8f/ILs62+60XYWMfjI35lijSQK8IYBJBm9O/XCrXsHuzkBAr6vRb4Jn7aLX
KvJHmBxlLNK5xsMi/iwsxckUapJHWUNFjQRbMS6/v5LtdHIq2x5VsPdFzlmyaR0M0pDowFCkRCEq
GGhx0+gYylFPJGefF0WcOdvNGm/6f/Ni0MGUBRc6DqKLQX51GPKS00xbaAJIpKaneRupiaQPhwMw
T3znYe3ODFCWmQiY5IkGx+vQuy4GO8lEHl9sv4TZgjJT4Ajo+2Ub8FOrxtV+zoNME+/iEzAzD4ZT
WOsZRhR2DwBPr7qMaRLI5JGboWOUc1d73A3G1sSmJFytL+BsXiOZ3ctC53duF6veOsnmFeYsMRS4
NMFVMZE2kN+w/90UBRCjkEpurbcPSLeiuBsDaJKp9qLnYl+KvOjSh1bMQFtcfGed6FnR5k/Mz/VT
LjwTI4ewFPxJ2qN2SnfMJKfbmYsK1Cv93ZNj/XcKV5dKa1tYx5nNHjypc1t/QXWCVm+LkujukXMc
ysUI8i8oflxP4J3RUPFhdKOPlbll1nTA0LOb1xmI+x1WYeKpBGnPpOVXRQPP91gPIMfwqfy8zRvc
7a7uSYw24YvkyLIjFdpQNVcmE0vk6Yamt6BYri1/ZJgispE4tQOK2nAiT3sGa/ANmrN8UPHO5IZP
KfNEz9xxsxfWKJ8HGZJttaBllVXJ0b3NpXbSioRNCp9ZkliYaAX1Epy6sLvSjAl+3Ug3yiIZOtC9
geSnMpHxnBZj+c6RdvTHe9BRTH/aEt2ePghBPPsLVHK/yJufDYWG1jrARzIBu+xqoD7K6A6gr4xy
u3btvgVyDJ0/4mCtJBxGXJSYSLgpLjj+46cfaYwcKhZ8Jx47alx5CWUAPOn3bA/Q2PwHlnWpztoo
NX3PfCex4UGfzaYk8iqNWtV2vtTf05zIfoFvt8gV7RUCuU4BxZsGYC0crHr0SuYMkYuhXdLZzpE5
KkgZ1NEjadnueoEbxTJ7pDhGm8+R1zx1txyZBiyv3EVDvycbTDyhA9jyOZ66FhW9j+Rv/h4XsLDF
03lupAp7XqUlfiGtEtTJM7LJ5ibpxP7QuG6fVwnO4ztci8cYi/vNY8yKGGWgJOoPqL6+3sfiTJHP
d0AV7T468sVZMAdNwDnVKUQKjSmWBXhXzBuiqKq/ajtuYw8stjicDBvmmoajIcWLpjuHNmT1TWMm
lAnmTSAJyFOSwikNuPU4c23EQGHxQCuNvqP/AinhpXS8ZwjySm2MunVTd2WqQ37DlCOfuuwYLhh+
WumvUg4c+M6kcZTyvABl6GDEp9WHUvf9R7Akfyuh2xotQfy3rE6w+EUX5dd9c1P9eqn+GDQCHd7L
e+lnNBoWNjemsX0yxw2GWcyfYMfe4vHhzsHi6C3WRpWSojHM5wBvCac+zH8Yojdo3ItAdd2NogaU
b6ig7aiz6UoEplgtIHUUtWerBH6pV5BgY9EEKeQsPlhKUQN1zvt9lZNsrEWJpYd2B+qdVsGB9pyM
fs70Ro9+Y0LOLmMIws/MCSxpxUqcBOEsmoJbgkf1dKh5StcYGtp07unk4W6/ZaEK/IY2i0jOj3yG
BjEWzQKgyQcRmV8+uVnUi305CNZ5JN/hqPm4/yBX1e1zbOx6HIQ3VPPirJwY2mJANiy0OhEgGjdl
dFyic08VqzRjDFRZB106M8bw/9jYBjomw8r4FyJt11iUozolJvOXayqsp3zKcU1H2smhPv/aZD1v
nhZfKrMF9yWmvPhQFvzeIgRMHIMDTaH6JZqgDU9Ka10uAzezKOOpc2AJtuYDlOUsARDqe7h/GUg0
JCkBLasH1qDMTmsQ+YLUKwQewZ3AWzUhvUqZENJzXMMFeMrzS1oF6NIr065Vlf9v9vOCxTvGvHkh
+PW4BfES229feJK1x8umLjYCkxcU+ugvRRxEAS0QgX9DIYkWxCyWYAPDjIGIEeZenmclKaoW9xMq
sk1gEpvyPalLK8/vfcgLktzp+X3vr+D2hUhWBFda8K4uffMw1lLLtsgvIzzrE5W0IajRQLDha+YM
q/DdQgb8JbDaHmNhZDlVzNKRaHPMK9fEsVG9bJEBsrRQ6ceTBeUYR3eyMa64lOAvr+X7phmVVR0i
R/jCm47zGrQJ5yqmOYD0hMfmruy4HpUVDA1GXCrpxQRmDFH5Wxf/xbhCAi3SplDV1Kf5o3PPXttu
JMBhH5wtDMzU0IfJAWTFKRK9NS0YvvLbaqMoA8zF5HZA0eg8QqMvJQ/xYETDMzDPX5eMV1zmYfhW
U/CfVkT0fWgK+qtblpUuf2S9tasLsQDtamb39n4bKyyw4lDwwXy7DIAaYF8ufEL30O8CaNoqCbHQ
3bsrwuqn3KBeK/f2P4y579lv5tW7NA28bHCUr1MyNrvKwrUrbmlwsrY4JjY/UxgWBbul1/iSjDRC
aJ5Bf4ut8MjHd+p/smaU88adnx7tjIClRXRZ1pV1qfVTQ+/Y2KoqIv8OFJnf1a6YAaIZAvV5wNQV
Qvv3lYgyPPZrAoyqCPGJU4QehjokB/BbA06A2wpKvAhCSd99bD752K5Hlz+TnYblejnMG7hEy2Fu
hCOopMh9b07PbAvYm6gOwFX8rPF1oUr1lzxxnI9ZLSb6Oc6OUW6+nLhUCvL5pGdz2Peu4e0efrmy
xk5k3bL2wDPC6kJa2wCNdZAcbVZqdFPyrHoji9yFcHdCbpXr8VuVrDWN8bb5TRnbw9domRj3L1JN
thO05THEo5Un24ik77oUUE2Z9phJappqrcKLn9s6T0c38gFvcqZl50B06OXvlaE37+WzdbUpNMeT
lVpUtgCRaEas6g/VhAN2+Df00/00CAf+1lbJVcV0VVNQmv4TYn8kIxIDYIj6tNG44MmT+CJTjae7
dte5HYz0GO4DkKjISx3W1lpzUfD+GdIdVM56hi3Ay262SZjSOySxzR6PswnVJd8Z+GqmfaPf0x/8
tUY/Rbf3Cm8zSsFaTS590NqonTy6EVkawgrJy4y22D4sJ/z6iN+eXQ+7ZOjSItqXtewEnX2o5wU6
5SCafVcNbqjKOsGGR3jYYpQDi18toDh8C8glGtO+RCqstUbibMZ5YVfWNx5XxW7eIYNu+84hBGpz
uliDRRe7FhpwMmhlahqIkrzP8JuACIYVAhDoy4Y14bTHPZLCmFBeTNeyT+U+tvcRL861KXFXeJCE
7wPPGjkn7X8C4MhG/hgwWvE/C8MUcFQzH4OZf2ypdvFuJsP/DhI4tmti67IFGNnAMoehYQQ+HRye
BNGrJg6wp4tMAtDRBS04+nFegf13WBAURWTKvBbWUsP/HpbD7e+vHMXR9mo/aCwNxLj2Nb0QCgsa
+QPzgaBwimpRDgD0qyhaVc1jmcygX1iCJgLQyPSNP4QYIqW+m9NNxmbFxdqKZjr3nhZvoe18mOLV
sLdqqbnPJJ4g+RSo2dT55iZR0E3VApPEqeqoK3ass93cv54qlNunUkJRrqPUrXwJVYdm7MkNorp5
/pVZM0rZ+N9vLsX9MZ/fMcJtSIIdRd9erDdyUZl7kTnx2XwxGZk6bgM+mXf6SXGinl1PKG0ngoe9
AnVkLBbZp9VrUSdtFAF1RsFmDZgZ/Kj9oYhVmtN+IG6EcGfhp8RWLwT3m3GgRcTXtB8GinWyPLjY
TFDLB4wn0iz81gq6QIArbCj5xJ0kSMuxoaV+UWRbRy3N3S6hi/WHyvyZCSGohOEgvo6/3jwQnTB8
I4Cvj3ufItCXw2R2PHe8dNvIBtgXPEjLeihVa4CK5CzR56TyAM6muWiM+wQDPCSB8nKEleDTp3kt
/zrN7wQspzZhnlIBClVs+huq0ldx6UhTKiA2OUKzlynC72GKlPayYKHFpXFSxNc4QifGwTmfE5LI
fxnkie10aNc1CaVSEd3xd6zfHKLAFDAuQE5bU+VavKbKzjHXKRrhYnb+E1u8HXASXspAptQLwZNZ
cHnB1p4YamxdJJe4tLVV30kiyVa/lKnRm8bKJOJqzNxBUArBss9yUOsmap9UWW0bB+JTxsatj6FN
+EYqtZSdV+YTMMOSit+XTb242KPmO2qrIJ2i5C7LaeqVusp9a9ONhoJP5cmJNtKufgoOnZlns48/
c9KVF4Ec6P1rHHtyT8tMemrOadie/KPpIC5zK/XDvMMuxlekdc3fddukOZgx/sanm2DnFqzLfAfb
Y3MbBXI2MEjtnd3LBJ3DJCb68q+6oUS3Y7JRyRNyuAVGeBUOVDqdhC3nvMHtEN5e8iAVj/uHH56q
1QFqqOJ8ckfFnRC0ykDMAclTqNbGqhziwTXJOS/XqP6/hZ8KhIKbySUdPfXvqeUG7sba1x7fpxOR
ACeACtr9lDYPsSfkvA0F7dhTDHtXHubtyilanolV0bDp8+4dOZp4E0fkkUL/3g9iYz0rJOJSAeRG
lYyO+WGReIXj1LdRE0owmcJ3EV+qp++opt0P3ddD7/K+w2sOm23d0EhiEvchly37XpkULwKD4k36
EmzyT80R/oY0N64cPh+XIdBLMT0DlNpu1MJKekvUgeFgsX8usM69zaIHJIX9hfuKer80O/8M11Z8
SMUIDDcHQtnlEO4pW2aUQz52cggUK+95vDP8LoZzJDqrwgdnKjQhtd2eSYdGrLb4ERRmkjUWxa3q
w2q+j4vAIuXHsuIqL5jqtnvpRj0tdsCeYxImCMWNNt861NmyoZD/KbZ2x/ydEpI5z3Q8k4gAxMMA
/xz4OZeUyCc28FZJ0wyVQlMzL/20ZzCAQ/OJidjqq67b1YMsauH6BVk+Y0aKecFKP7H2k1ln+TP1
IYhiVW99qs5McJ4WKtunxMlHf4/MnQGmZJNmiOzC0/+ewa5Lvr0GIwE2RrLK4lcPmJbfaZ77CzMq
X7pVV+ile/RWTrd04In2psVsy9u02gJ9yLX7bhzua1iiIa8VhDdRET39sqoT5kCtU0hMExLImcHk
Jz5s2o7bT52pfcvcUDDEJ1oLDrvkOsTBlxS/ZyyUPQRNQ507MQQ39i4dQgJARxZNkUMwUotL+BmR
tkLlXW/ORg7P+fGAQ0em58/q56CepxHqlOKitWzyseoI0rVYwP6y4SqNx7NFLYNiMbNSA9ezCK+m
bKcepyAfWWnmbL7zE7yMeMv+vi6U6mPFWXIojO7rNTcjkK7UmXXdtlmEvXCfGaQW8ys6Nmh/IxGz
EAN87Z9MInm77ZJJwEhJ9KJpCs+BqAcQVttVL+9/SAjsuuQYoBZfc9+NivA1or7bIryViDXJMm8X
TGGcE4iLbkN6Rxn8S8fmOSciUY7WCDi6TcwLM0CKatkKS9BtJa03GQ6yDYAiz38q7pYHfrsRavp4
VPCouPcaCiMXmyM5sMjyl9Ic9jp9B3dDxvftf8v4mVLIxOiCAl8hxR6U4FHEagNdXwxHMCJUE6ts
Goxlf0UyTzA5tdrxTo3ZEtA3kiGnUp+nC6EfrP0bsUiCIrQ2geU8gMkMyLa8ex8UbqeCnHiRKO3v
RFzg7N0IZv+A1bmd40Oba6VOOwqMMM7HhfjAOXFjlzN9sYuz+0GYOjssCbC7b9CQR6+dKuXTasbi
wb6EGzCE4gCil/LYqyOMozyiQD5cpkUQDLeASB8R+hBAEdE4M5KaFbyLPDvpNItPWSrwjc0B7efq
r8e6SrZ/5BvMq/IsrlD9P29Zow4mmWmndwtO2UDFSOl9sZn2XjAxHACcRh7rveX7pFmifKoqfSYI
sCJO5mrMAu+Y1L+PWmpiHqsC2SEQga0cfyvBwKFq0xzM8sh0+17Gnkm5bu/eAY1H5dd61CbrWcIx
d+1hgBElOC6B2JFj5vtHT5lzq0dc19Su6EysPCQDopUujNMkQR7u3IEibzyQzMHZd5C8rircK9k+
5tYPnD8s/Rleu/qYPl0XH/NoQnxTxdQdavgF4spMOJ++SY5Dz8oOY+0zuHZdvGMN774l6y2WTHHS
G9sZSfPsJVYKp5c0xQwq0GpyzK1avuuNKikTi//tt3sZUIypcTTDlCeAGfUt9ryOaQRjkBAf7PQr
yhR4X+VAYETSpRZEmC3hcHxP8lRHlkEourM5vix8Fx7NaF4tYrgYKWjyFx9MyetxP4DuneSKFdO5
10J0oL16HMQrpBEK2I/p07izBeeA/tR3EEFNVyvwzqd5ceqnrEanmpMhVwXIaG9drkZwRRIMoHs7
EmAppy6ybVeXrjr9hqrUJM0zmhAjbV1onAGURSgWi3z8GHtvEQTN8VHsOdK4Qv6rjrfoY5dARGgj
5U8wXM4Td59hrv1TdkOOOH7JIu121sfi98wc20/tqc0QFPU2qupE2hreqot4f/A23+r/4UvmSJTF
fTMseF9WXURZMzEUclbVvBVpynZhE0Bm9JELnmNOMP4hCgPr8jDYER2xaFNE3RyReEA2TdqEb31F
DbAxBY7qA6QT8Fc89xMp04nuOQmGFaZWD2NmLjv0GNqFLD36rXwQ0E7rbtR45Oa4pgEWH70iAHYR
r128lNT+Epr/SLOEMVdZ3vIWIyTWAYzJ4oOphx7Xy1PygEMLkzZSxZpIIVjKvSS4v7xL1C706FUP
Aoct9dRs6cjAfNXy+1zK76SYDTsFpajyQW8IIFHjOG9k50YB/2yRRIjY9pTgkYdZH7HcNnKz9rFm
PFto3251+TMXeDQcRaDAkGdj3Q9scc5ItJUaTQqINh57tqE7VNyAiFXK8lazSvJ3D0KV7s8h0Y1k
hwPkSotmNPoGVQENyRB3ZeGOmrKbrByomFbWYbLt3lsBQ8XR3UYig2EEpKKRNwyoKS6Z21efu58j
kNrNyqxlo2sV0cGULfE7zYipIzb10kM7XWsl9jwxTlj6KxMt+7ZX5Tm5AcYJSvFRNGyqNUlwNGTx
ni6juqeq2NDv6n4TBIwR89XZ7/Ex9vjmCYewM97P6didvbhpRPAnIIqUuyevx0S1dKVsY26lp8W1
7PGug3YQJbNAq6OsJbb97bURzzavkc6Y4OyOSEfSY1GKSkXOpEdwiMuGhUmu8Fte/zBFWegZMhRp
4cHziV/HQP20MSr+iKqgWo38M+8SuWHlxliDd0GwX4cGia2SuJIEcLzwHhvZeUOP81p/ENMs9lKi
GFb3RSj1XEvPQfLAKneaz5AeVk87ys3MYZd/TH8UBAoSODyt0iJqBeZTT/R/VRlL6fpEzaM+dk9D
AL98RiNqLyEPHV240HkAVD2vYz8TVPr68qhFGzO+iipoUgtP0wUjHni6QV8d9KZrgAoept9C7C9R
OykV0ZUc31Aax9YxF+taze6mvBUBernk0mE4sRaadrplfHbnGXU/8O5H/UC7+Wsaoj7b4jv4osAT
ckoPWDcJzfcXgpTkO0S1XqCAM1RogY85aYdtsNNghMzMBj8bm06Ox9x2hrIfBhXFkFAALnmyI+7q
krUIG1NKMVr8ABXASXtPDX5YNmnoVXxQViyW750jSaUzYCjTRAObnoRtnZJi6JfVzH23cAQKEnWZ
Brtdmch4EZJLNLKk5VRVuSWD2XOcZ+0tzHBeacIMhUgUBdt2f07CRzTvJCDFZEVVWATGGSdIl6tg
Eon35IewnXk4pSMZwJAwiRsq+E8ifA47rz/KLqwgGKSeRyowpvxhwgQDPqwuD47meBwXKnILcAQQ
jzSmkG5Pb7vwICw/eeWZ2dhQIzV2Gj/MIsZHrzXuEKgYiJ3HgcmauaRTcfNJ2xLwdH5GJVy4tWCK
yy9cRBGAcRafFdJNyEeuPgZeAsDBNe3c1Ra2lhBsoAt3jPB0tMty+AdynswTogFLLxi0GTgc/1HP
Ef6jJV7yOMWkQqmZH3MkwUb2wLdc4BjUhof7oJUtbhXBd2775eBDmMjcLGdUQ5lnWt3CeSe8vvzy
BI0Cm+lsQEikTtSoiHjQOx6VIlcNLKB1TbVS4s4xx3Q8XbigsLYFV+Hf32VoiE2fKnnrRRLxrRYL
OE/QMRwNCl7op4LnE4wiADSu3vSGkZUPgXTJgfCkCIXcw2AAWgaFup/+8dX3OqIwqNfdVkGvS7EH
CRd9aWyw0N8n1rlRpfxn9Hz8zUg4JyVDzVGxExU261TyF6/ZuFA8rZQKTevG4q6+fXJV8/qzgkr/
6HE1ygZSYB/qhwRVe195Y3vOt+8GqazQhy+Tt5Uwuj4hYjwkSWg5oEVAuQtO/IpmZt2zNefAa2Rz
Vzu41r+KH+P+I8hUb60QC+80P5bLmoVVN8hbzaAcp7aSk0A1e/s0dQdcQoephUD2o1MginWHz7Uy
MxJ1e252UCKjGLWCsJ43ZB98OIaMnwe9J0nTU7/JTBmjT/BmzJ3OXEPvqHM5hBY4ZxZSLqpobEx7
wTv82i0HznYSjBrnMX3NGzxQCO1sFxssJv8FBE3BRCdU8k1VBtn0FawJ6yyzpOnn/asxAz4mkeeu
dVqKFi39LVZsY9XsZ5Ve6TdvA4fyh418x5U35vHxKp0brIgoCgnFAb9xRCnIpzxMRa5iZMmSzye5
h8swhgHOfgg32B/+Yz8RfFVAas7UICkbNafqoXEsISjgv+zQXN1Gz1X6PhUTtlEyoYRY1XnNs8e5
LnNAEHwVO3JifLcGZyvc2Gq9Gl/S76VGPALRmQLJm5h1ciRJwXgQvGv0AjtC92QPtHAkK3Q0RMpX
SrnnRlnyuh5XVdGd9q0Rokavbk4Wo3d5EomCE3iWjW7TfvwHG8Ib8bgCvTSt3VdQz5ZekzGjqZ+q
NE8htb9J/kSQ0XUy9I8yl2z7q3OKwhYJ3bwJYJSe0u4BQJr0PqWgK4i+HJJARLOvJlEbgb3+8yE1
TlP/temJ0Y+LPAjrLrHeQMOK6SgidGla90C94vQb4KyS+6ZLB5aAW8ZH2nizlzB97wHGLKlcpFnH
tQDn3XXhX9ZDaV75Lmx64EP02aPzMIvMNcbyN7n9jwAy/JEPjCIqdTNjOGUq/1d5NjBH7i5vSa5W
q1biYqRfcMrzaX+qFaMVnO/cErs5HibpSpLYplsZ6ZpQYBu4k02YMv0kj4HiNmJcPNVOPRKc7eI5
IeS4dSOQqYP70Wtqh7JpX6nK4aWXEsvjdWej3Q/B3oUShbwYapImuWqSHx1lElr62mIvcBrTEBO6
Cvtikt+tz4+XFVXg+FKsQjDnUN+W/6v2+MYfGdZ1ZI9YEhwgijX7lr6OTAh64E4C69Mwn9BBpaRi
uJjFRKja9K/wdgI49wWt/MAMMPsqZEA+UA1bCepQHtuiNuyCMfKqJfeMY1YOU+ixD8mOkkOsoI3Q
ExmrnEhlgTfRDNe6CrahlcGSipiX3Hy3bhLUo97v8Y6gYaYM1GDqouafWSkMMbAbggEsZYUskeTj
LbH3cP4jZJ7j0gb2e6+trL7bBwjcpj23pOh0OdFD6eXgs8eT23F3nssvVxrZTKp1rm5m4kyQdJCi
sjnV7771EIopb3pLBD5++Qgw0WHWfnl3BqBoLkp6wCsV+aumOIQBh3XjEZKfcxnwJEfsu+iiowJU
dVtzFr9tUIUXesKbHRZP5Z3uLy92jDIdoFK12I2QQ9Cj2JxV61X/kVUd36ok7wFWny6l+MI80BUg
VjrgtubZt232O6F5WcRAndp+E6enYuIka+EqHJDBLAZPPS6FvXP5rKjxJkGdq4ImoIT5xi26exVx
IUj2MQPKyEhkMD6Fwbgzk1OMRcovyWcOQbxEjSqyUtJVO+7rD2Fgcg8BhZruxoVuPi+IXYhHg/49
D9hp8PjcEmtK6dM1MYbZwwDXOnpKIYGEAf8W9va9emHHzjBtz5aH2AVmiSrBijbOPJlh40iPpTz/
GL3dkjoJ//rt4ecMykGdUttgZWCHbzUl3pUySC0pKS5DsKavc7X5wOMxtyAiaxlXCzEO6bD53zCI
fg91dJzq1VMYtH9BgoFv/A7z14b22SNQJhIKKP2qfNRXMuyuwkzdM/L+1sT5FfkV0+oXmbXbJH8s
I3M+Cb/o0fLLwh+4g0RfOSQ7iVizps0EkhOkgdt2+t9yW53QNg5JkfGXApGGGr3ZxcjngPBX633d
MGi2b4cqLUFfMwZuzqVqOEoXQPzc79rdAPejMYIG5haKNfIP31/WKRhIeG/kdptUIAioqZ38v4FC
8KnSMnfneIW8lQJa6lowv4CZEjzEXy0nxrftuR140IRYuVAWmjsIHn7IczRDaSZckqPszSoexNVx
zW3/AvMeJC5kGNzPbzduib7BFkKMFoXTWQd+2/nySFy4OWYaZm3e/3PM/GzpHrjNHjZ6WrJzhv6C
EKuQmqSkTdMCtQjlpO3+edB2MAsen5bozJFAlIKpgoK9JIZFOuwPQU3vAH9a9xvGYUg/eJqjDgTP
XdOPKV5MgUtpwoH9zvh8xxPq/Zrkq+MJTbHfe0H2VW3R2auUzP2DlkVem/EKOiZ3BKWxZcZqowvp
aOVDynAaonTwE2ZjT7ccWwFpWlijlqd1OuK7Nk7l1GhhtPT0lVlqXMZS//3zRN2/eCWD3rZjBZm/
5CunX/AxkalMkrhiwu/m0KSza2Js+jWNot4H+ux2GEOEs3+tiMaGdpNPoshj/54JAQUA6rID7H18
e1G6uZCweHbBu4aaMN6artX6uGNctTW8Y5eEAZODCpJkWEB7XSYwX7mL4WyiL0IhqQJOwsdnisSt
wk1RvTj4NXNjKhh2dgrHrQfyFNdow+XO4Kb15VvnzrGfyoxx+KwjgjkQs51EFfLU4nZTwn9LCj+7
1xBJ3H6KIdvMZ4bCSXeYHBU1uRrhOIRKLHJqVPM/ObPxMSvuhSfsVhlg8MMXQrWGrZQkX1HA8Y7Q
ZfExzEN9eQB59L01z4o28j90/JqP8UzffECyzHS0R5gC1NfKDu8mLq5ydEzuMQgNsnbn6nPpSIi8
NzVUOdz35oLb4d+7qLJ8dTs4JFjxPHxrxbUmjmo7T6oFWoGUHU+6ZBFgJBEaDTZtjhQd8Cyl928i
NlFM0He8JdbR3aXTX4WKk9LXZwipwYil6F9N/gEa+T++J+tF1YfTXHH/FGU+OT+0KbLQjIAoDxIp
m7u97GoKhYZcdRMpNzFGBR+P3RhVG1xJmZBQwxdos1fIbZIqT1046LpgSzUGhOrf7a0ytjrynpnh
y/DwqR5V+ffr4Hm5mXD109tUbYnL3Rj1Y3nUcHy+Ep4JxOhWO0m5j0u0e1MsNDdNzdBie77cLQIT
AgFavvJojUHlzwGZEeLL2B1iCY4+ldgghHg5ZWYotSObrsK/SKeQydZFQXMnf6c75n+yAYkUn7zd
8iGzkrx1jq1pvON8ut/p1vVGS1p88kn/cK+Ex/XiVW29JPgcyDKauKfCcoAJO0Z/rKsX/jb9kwP2
SHYxx6kpP1TS/zHrzNWGGQqOV3EFZV120oJgG0dlOZ7j5/3rXONifaU+PMFzlmw+I7zaO6X1ajpz
zLibeXf1LlV6rE/6B3MLaO+EfO8SPGh2VtFXNr941wkIVeaAPGy+jbNoBYhmPB0Yxf2/4M/UF94Q
aINV3jDJJdGOjJOfQZBeuV8t4/O0xKPNfF0WOknmNoeiVf0/ZZoYeAiH4oezbzoWpH9vO9R0o5AZ
K5b+9xU8iCoXNOgoUawsUAC8XlUaOVYCk3RZcnKj6I/8POlAubY+wghquoGWqqwdZ2yuyTeZYkUR
D/Cwk9W7ljQ7hDo8qI8TBgZrsp4fvzCMJX7HgHivZjJ2Oa9YUx+Zk1xBLILYpMBf8Em6eA6k/xql
Wa03V+Vf+c9syUU7plO2kUxCC5HvQzWoSV4mL6CzchbfUwvyf13XFS6/uwKVu+KAUzq99oMntpEN
HkyOioztqr5Wf29/QGFuR6Imsanx9echSk19i43Jnt2CIe+zVHzrDtexwvd+cKabOh/k9IkN7gsU
TzGou9O7t5yjuWqopAYiZMXhWD1qWa+eXHJbKPUkT8zP6l/nhCLWfDcxUk8NtcevSw02k9brmfHJ
nsbGV33ibxymh2uDB6HswZWni0wBJwdmTOf+XgvKKU8p/pe4YH3EHDmasndacV3Ia6sZiGNeAFkU
fK9WTIugCOdzvvUZiXVzqutJQ4xDVZa/yyQ0Mx74ppqDQi63PUpLjEQwMkAJS30LWJXXwcvRu8Qt
kKiqkAwDaTFrVAp7SNuYETKGsF1CYCQ5XYq8SQNwxswZvY37h0xm75ub4IQK009vhx1Jnyeh5+MQ
rci0236oNBh71wlseb/9si1k8b7jFFn6i0djwQ/IYw+bKPWwCwVbwA3ytLPbG/jtlXAgmR/x7HYH
kpiuLTPEycQH0zTS0X7frCW1Kjpx4bZGGLxE2bKgG7A1OzXIIT94JDo7ypAzM39/YqqfinxQ0SaX
+5Uyl4j0WSy3JHWyCosEKWu+Pala7YN9KADGQuSJCHx513YV3LKKN1IwL0ECU2hE0HTA0147VUjC
D5ZvYgOK5htz7dAmosslU5TMhg/TMLAfeZVYHlC0DOg1gjK8NF+O+XKLq8sW/748s1kt6zODsY6W
39rcojhV9do+kuLk+yrZnX+bBtn74NVP7hsbff3xNnfhF3X6C/dRQk9MVck6VJPVKyeNIH77jRuv
sPqOGgTi8QI02AtzBO8pxyRx4dJ2xrVFsJ1BSJfw2KhwkQzw0IkoSQtF2MVhl1RvYE8BHgiDDeX7
RNp6ur8RsO8Z4Rf5n3Bf9Y8yNWONB4qkTFDehm9u1uQr8Q8IOplxjfdPs6GE9XCWOG171ChDYHUB
ymjBVb+6h50WDZFpetLlxa9BhshIxrhyVVN7cLaHKHVjIwarMM5guok+uFuTpIgfe3Bm64NgGDhD
KEpHQY+8Ml3rQHm8YcGwTzsKOCH979WkVlepakVkbKor/vi47Zv7SLF9nYQHsFpnIqAaFX5qg/A2
LN0y6kf87QUWLY5QJW6Y5KLvuXrtyhYfgMBrgf1jgWN9srfhGpbPVL3Ut7skn47hE6AhO0o8NT55
rZwV7HRX8Bpr+Y2mD5ARsMsJdlh0L+3QQTHiv5QsikqZJ2y7+a6wRsLYoPA5RqvZulTdMYUURGOb
lWJJ6mnEt1hW5PHHPjKtf13lhasiYLVbawJzgD9mjTxKqr+EjAkmfIq3lG/yyT+iPeuo2+a7dnYz
LD8JbGs+rOjSU1CeW9+Bw1keOMNBpAulxwloJ5owCd3L6GzbtGxVOmnS57HnYi0QzLzUTL0dOWtK
fJTvHsuwSR3YHsVN4cPG4Ghwk2zGUeBRwVXoqVgnYEdldAd2jUN2rdYF/SRCbAZvS4IY05IDLoae
vCsbaPHnBArw3P3ckIzc2ZCrmWH1jUknk/JBwFtYqX2u6y9wZPuZRz9u0828FhiAn1V0m+gfpe99
MZyGTkh9OQLL8mguvaSHv+mwTZEqvkobMc3oEeUAtk6ZuZc6g7efuWeC7xc98zzbhLsilq0BQWFw
qdActC7RJ2fsTd1OC9iM2s/cps17wjpZoBGqGmA+Svy9thjCuvrPoz7BOo/oUYqo4EZltuhIUEju
aMxTaduTMf7o8VkwNUg6mZRR2SFCEz8MxVs41GzytS6iBoO4RcHCUPltvFk4m6dD3JOoEIq2WbeC
FDpqWlr9JdHYA1pQsLxhalUWXt/XiCxvSz8//kgBS413oeYb6hmLeweJZCOzoUMg6h4d+EOTfkHS
pyhezmFlOvVWg4VqdK0BbDS3HH2iTfUK6Gd/+8AsBghcF7LaXyFFCiIiEyMlcB4ogPStnzHt9br4
IvoqzeYOxoXKSuYc+WvAw0mwVS11MlNdrCzLQTMPqYQ0GSLGhaqpG6ESoT8DlCvCBiD/YQyyb8FF
tmFZMOTquHNu5FOBt0iyyogmvW8gVhT874Fht27U2v9FljVyJDoxjqFJYcoCihYxk2RuiSRym8Gy
jzeUqV2W7rh6I/2LgxSScxU92m8KLgfS2/Tpe6otDaAiYbBP1NjxrlJ+Ye4xHIG82gk32ihOkHsa
SqvvAKiO+YP3Wsa25Yq6GuhGvUqjaD13cM0FpaYQ3NHwGXj/nyzWJnqYl3taD9GnRl9Jjm5Mgf5g
B0Uk8iELxibJW7PwR9M/12Vv7NJsg0lQF72gXX7FtxrcUeImv13sWSESDztSkaz1bCrCaCDHbO7J
Lm7Pl9LfKfDvOHItQVAZxe+/2AGhA7ye1txyU59i4PVJtskmUt1nIqEnI1lmJ2t0+HE76xMcgepC
jM+cLz7NvPy8p+M/nevCRdlJLMBzD7jaHbihWvhbe5kao1dLvn5fBG86Aup5EiZ2CUHZTncJvqQ1
LHuePGIsB7fw2oNBB8I6N7TQ8rvGI6MAs0Iqw4HodcKeZEI1jK7pJyv9WWi01gtjclBmMoZNEBG5
TRCYapLX9wXHBbkvIp8rC6+TFpDvu1/yZxqjSmXZWv5o6V+PpYtHxQl0qWA3ZvEE96UF8PSXl+/w
e0KILSd20zeEwsR493GrQfAlznq3BihgNH/qlRauwmL/4q4dCYmeoUoBIiZmPle4izg14hAL5Gun
miIhobwi9u/d0CLe4QP0qU20wO0OsFunukrEYTpx1/fKwUDbOzm0c1Pj4Tb/HxgM96PQNycQbqrA
gyzfzyqyFO5LbBl6U7Mx64wWi1TvebBpWPLKX/XophRFPx9n2I3Z+QH0UxM6Xn4N9p+fTilHzNow
x02O0DTBbigrbZRfQLgjgEWbnYVbeIaJQBz5ulO821+fV3AFM6s5mNh4D3I/irtJa7LKRDbbM2Of
QIma7yYvHRdT/iPJk9PZhAyJtOdRTXeALYfYcaxdl1os9z3O+ctlc8KsGEookc06YzBi+mifRo+w
gAKQBlF1x8Tr1yhONYH+5rT0RL7QOBluhYe2JcpxL0kI9FF6pzJui51z8+KFfGxgXIkElNY7vPzd
NEdH6Pxp79wDDWhbsSIGa/AEdFfFnEpgvB1+hz3AtxVMrGf6t3bl6IluXTL05NfgMt9vVRQEDr07
BGDNySZX+lliTOUlO7SFXbXAX0zwO7E2ptr2ZTMJepdWR1KSPhfHD5s=
`protect end_protected
