-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tG0dyzrkktQ8/86ZUf+HTw1FL5QvQhEv+IDHR4mdG847PhoMhDXhuD/K+Inu+LejOLWpBWV/uX6E
4UvezwUUpWnL2bK1p+A3JPNstYJu6g5BebiFyjYJeO36yRrm+xlL8dWb/5fjTh0m1KwsLvtGHMBY
LiRFgdra1jJ4EoZW2sI0mieh6KQXIG5fWnna339/vM1G+JqrAvPF7Xvj+1OzzMCo8G86o0oSopej
0+ERJl6g240mY0VVypdBEKUF2w1/JCkYHFzlv9ddqHViNUOlgVG2Mmk3PIdFP9oL4+qxucjNiMRb
q3Ng8PWaEmmwMNQWgvDiIdJcFJq/o/arayiGPQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 22000)
`protect data_block
D/nWIzhme8XI8FCT4RafLZWpfFWZEHHa2iRbSM4MdfgA3NoR3ZVnFJH6vTrpCz8886VKHyfzd7IX
qhDSDWmJhso020V26mnPkiBG5iWXqChKuSbGj8x6wRbebAdoFctc8Z0fzqNY/RZItqI2WvKi63uN
gjqnuv06bLq+0aWDCOgR+TqoPZ9viIu0kfALJMu9OKXS1NqZTPuRuuFg8b8D5DG1aGfvJJGR3cEd
0Xrb5zfyAHVXBrbOarLbdv6uC3KwVM9isYTFFO/PuYQk5jjYKkYW+EfEYTd0JrusV56LgMngz/Aj
Gqohk+MsvYMJivF6yx94wA5p+0VvvplVEeTv9oRT/1eZX0UZihC0n+Hq3T5j9y1JmvTTkg+Jzpwv
lnSOGNweDTBaNGQ0CIiUFLQ3/be2fZocmghFrKEbSEqUPRk5vXkc0MNwUMfSsC3UOW7tdx7SVFFH
nAZ5dM8kF7epPtgBVeCbEjVUzYb6M+uUokhAXEcNsDhtulHLQv+ekR7cpZ3akU/8CElZuK1p1T4A
/SgLRGAFPPFEko8ZSe26PNDdVtCs8OSMKhrRh9xsT9DB/u6hi8S78OuOwFHcD++6VD7SqyRMWz3o
n2ZeCyfzTUoWC93TSGNkRXrazp3/46zyPIh8PtblRsCtIkcvzbNRRmdkd0+tZ75gWJQnGMdms5a3
w9QAGZcIPUx7dlvwBMzvajmXbAUUR7gmrODGF+6dhaRSFwy/IMkc0bikgkCH9j06eVCaaMZPgYbh
HlrXyDQBN3Ob6i28+Yv6bMEtZe7muitPGIWJASVRbfuHsnlc8kVnbwluBJ3exC5I4DzhMf0AdMaw
QG5GzRkPHaNd9Bfld9wYwV2NpAREVPO9I5Xdquxk1qhlH+3StAerTQMEDPOS1J4lRupRsq4TjQCe
sOtUjajqVs99PSWylBcIuSzvvHsmbxMoL/XL6x4CRpUhrceF3hahxfAaf1lDjQfjFrLnS/6BWFNv
0OHjmuYOEVi8+MD6GFtGb5vkm4mue/8omlO5QL+Mx272CwfoyYpR6cdOGv0SJ6i9wYbPme9Gakzl
k86sF4P402yzW9/SGYanvH9VUD5qzwBvW0FsjxnwYOgNjljShwg+RuzZ5Gp8K86Dp9alqAgPbfL6
jG79akgVdmgOyFwRaGfzRvy+GLBG3p+0lbUW1I2eTx8VTQ/juCHSUfRl0vMr3tIxe6MPD9EXC3Gk
oEtXw7tTk6TLYHPImQyUQVje7k5NoTs3uUeMJ6HVDW8SaI3Wj/PWDNVYlFsDX6ZAQ/NeAPsD3FaV
i0vUek3D0kh9yjUj1LwSvDoVep0jRQAfiLq/5izl1Cfg/6gmpDgf0ixxk4fn2LE9BQOZ+Ovkx7Jn
PT6si4AlWEPhXYH+MnDLpqS4+8yeJWp0SfQZp1jLG9E/h8mkNWnTWpH2Jm8CTg+cmd/dfZDtdXvF
NBMhttxUCehYzB6ztavAl/YJU+HM4kf8swS6qNIr05iF4z0AGqCcuCyTIs/swJIOIhK/VPa5NpXq
JsqhYWwuY8oWMoFD5enewNnL/vTiEC3itMFBK7lsT3HGT1s3jwU4h+EBWZCsFDT2RWXlQ3MDBe32
/fL9/dALPwB9pdigY3DevBZ0GLGDDMg6BV97noLZ4IwNZTVvq3SU7tqgye0yng3Ud4fs3mq5f199
elbbTJiYAXt83F6yqiUC2uYCG5aZALMcTEHj4QBHsJ5FjI9jKWBgw862hbf1lad0zhaD+cU4xA5G
UdoNw58XUxF10AO0oelH7t3syLwZ/K9BCVhlRUej00VBSsZedjN0VPHNiQ11VqVnJgssaL0ydusU
CrR9Dl2pf3K9ODBk3h0fOYjA8izqkNsuegcshrIu5Hpq+Slk0BZ1rtuWVV8OiQRqmHR6/D2ST99N
Sfc7yw7YJKa9N6KOG5/DstwrZhHBnHHTCZ2LsmJ19HiL/T0xhdJnq3upXzQ3QteGCGXbSjnkq6yC
ZQTZXlXZrIEemsfO2PsGqJjcE4Cm+h5/PnIVoO0YmenThKj+lT4AbBzQOQ+YNH+awkJtaMmZVzzt
ULvDwpjygeyS0b5RPrjIOQWrfWU+lp4qRso0YRYjpjJ3HV27gkNjt/W9uTSyiBlrYhLJWCn358sT
fy1I0BzM1nYt22n/X3pF7TWtK2VCf19a66Lb/u1HMUPpoVJ3rcLmRE3fkhPb3tcK1zWC2rUcksvJ
ZLpbmNlf635NGN1N87FoO5b9cVTQe9xVyNbPzCrUSUB4h4BgxaYBhFUpfiXEKecdkJBSyicm637X
dtKtFxgmT6Lu0irNp2J0x13ZKeH6en9yZReJXoED/7mZYkUuGQ0i6+2rfv0VXURzgNxALZR6ZjDn
gpUY296FXFnh4SnW3xrYE/9bYdkMIMy+glhoYFF8GfeSHtKlUj/arB96qSdFNVGwNcqM/30LxPpi
oiHsArGMUTwMf6cJw2/38dWLW9c05vAT+dNIZkwFBOclQitb0es+cq7GgLAIsxcPHfojehdx4izy
YWCgapJxl8CMhdg3V624B67ZXbLhmNQHXQZtIDH8EKbymtG2iCAMbNNJ1QP1tBi1g1+ubAjWtWzv
LImSJjkOX4nP5Hjpis2fTtC+Mf51basziwx5p5o7wudb7Mm1O9birWT4r6AkHvFDEhB5PnVafYn5
Sox1YB5zRTO461mNmVkRSFw26Kw4tOAxI3GvkSV5cxe7NWWmgPURDklsErV2qefz5Fqfp9aMk21N
mMJ0FkmGidJ+LX73oAvARKMqee/3o1F9/vLFez+0GysZ7lkKX+IRBWlKM9J3Ilj9Qv+98AHRR8d9
BeW1FmUSR9VMcrUFxf8T/Oj92R/QEEwbrUmNNCiz2m+owussUczLh+jv/ADN4mKPdhufGlJhRK7X
rKrUbur8Dz6TlVXX5eiUlL9poATZkfohAiIquirYheuStIZqaLFhN7KYve4PxAPRadQmrEpX1TNt
HGFzj+Vqk42l0eTVsF2Y/3AQ0mUxcsjclDVilfA+nfgmLv9okGN3kIb7z7iznc3dNnMjPjpMw0OF
Y3D23vvWG3d/vO81Qrt6mx9qJwDRDTLkcau5g6Ndai0sx3dG6zCFvU5rfi+KAIkHhd8av4COEjuT
9Hrb9gGWTYOaHJ/Ag7tNg2y5YiwEDOs2MoN6U5RS7FRQDwHnpiTkqPswSPWRVhXadFYQjIKkhRdR
W76eYc4DobevQA5vSbCVWdwIqZu+BsXZXgXncYPgb8voSfJhgGro5WFGK5i2g6tQtVpJkK/PT79r
f6KPow05UPjj936d9oCZpyYXcf3QkorSM114tBSlJnre1NISGkrvieMh7zS5DTNg9Bnn735awxMX
Qow9JI4PnLFDjPjrWNNT7lUWPaoc8n4HWOOwMppjYXRsmGrrFZ1dXQ5Ew+cPBJIitL/Qj3LeSJYj
ludjwkLi5RRm3PRColpG5Nj9fYRF0YqVzSDE5u/XqxJnfyGKNiDwoFiSng3m7GNF+bT0PVQTdXzj
5MUc3Ewp7g+PI4yynmfA/ByY4LmiaQDRne9EaFruzwGobHIqWzGw7oEF+NyN9AaLEu7cXcT4I+QS
Sz0wtPEmKwh5Bm0HA6E/GnGvLECNEB6v67pd9EVJYXdJyk4PXFgupxEYzNUaNy2045LKjgw0rEQf
GiED+Oife7HDxoqVRo7nyTZfn0Lfg4fbtM+jh0Og5s7JE5tD3JRu2RyE7RXHwqaKfRqubNUnRk5q
ztx3+t88HxFSanXTVTNuxE3iGCMBU3n3jHqf7PFLMduQ80SlRSmc9fckk0vDtgkg6qGfTSi/ayQY
kjev2AbUxAOS3KSb+UYqPSNPkMkQnAiDxNfrN+nnPK2QBOk0FHKUBLhGtvY5SzzaUr0rSsee6f7M
okHroaBJACFrDaE6dLD9VnVdW1LIEd3VVnflEouRT1kvax4+eIpMHVOQ25YyyFSWRstqSHQpL8e3
alG8f5S45IocTIB4b1Zaa1dkPPwjZ5iV70oxClzC6/708Ie3YXPs8fXR4EVsTy5SVCD/2zzcdxOG
k3iiKagiGLBs2fnm/SLUNy4pblDDRUXsc152sil36Kt8C/5kH5McpeOh/M31AyQgFEKAifqcGL62
cgmhOkJXUVtbb8j34OZ+pg6o2M1TbkNXuOs6OhaHhHOrNCObATDYMK0YMh9jZs4v3ywqqGA/ueqI
nwOCkO3Ud49/0rVTv57SIJ13ejD3HyypGC/5W0GVwwWLe3QEdjLGpO9HBjIUM4WjjZVHW7q4Po0N
l7KD/6AoX/2BqY3nfV1KejNL49G9iraA0srA9UzH7LrchgiXHXjt9SIkxqnkR/jMyikqRuExbzYX
G8L2gaOvvOtH9C0tVpM2/OnFbwDFEmAjTXbkM6jdN4YvQJulLoqRTqBN7fMlZfE8jsXCkOCTI54Y
zLZL3/RANS/tWT9V686WhzA+LLr/4WGzPTnZ4TR1Fq4KZZzuOfx8PU+ZbIjz70RRACOKclJ6FCq9
PJO+PLQjtHXL3WqgVrsUTsNtqVzT2JLJOUyy5YNLl8cvgwTsav9BmhxE5EPrqjug0hhn9uBtfuWM
GDFbsYLktADEZJ+SuBHqPPfwJZe7wuUcCSGOfR0bD+6bfnkSq4RfJHxB5qoRe16CTtgPL/Z0z2vu
Rvdbynf8MB1yQYzZUG1F0NthMVxgOZs8G1Al8mhy0CkshKkCnZZMeQxvlxT9Vc9t8YpJcY+XSO/4
UXaiqjSxv5pr3AItFMFF+hcjAwK3sBeIfALlg4XV66GwcNCLfVIZhk98JwIWLybOoC7M8k4wANwC
71PVvMPCENiQxgaRrsItXuvB9DojAGZjwGtrhrdPZJKWOOOhMF/YgpOM4ACToiQDreOtk3fzThQE
qwfzhtqr/ulMgv6wkla6bowRcF4lOIJYqGCY03DOlHu8hA26BImPzpF9Uur16fA9/6Rjg+v7qPXZ
DnzXRSBue3/lKhGYjL5y/X6nFleizCk50jp2DIvv+9vdEcULsXBdfwO7uJgLjvwbZAa/q6/akIml
iCyjGyoI2WjxEROEIC/Tj40bViQRXIFwRUFyzcoL8Zyl98b3V57dAWRPa6zRw89mVxQbnpA+zxHo
r6sbXhaMzE7o/XqUenvK7uq53XAZ3JaXScgBDy2+RTI52MfgRvtmvohbFyMvwfN5N92Zlz65haEp
bFAisBytb83wn8qtf7b0u4CRvEEoJ2jeAxqit7rp4l6vEyMAlkbSJQare+Yv6+x+Q9AdkP13ZJFw
umNExlQ9kC8AInahEF0vWV1iMmDb2aqrks9/ESpKnM28vXxKpivJHIPpqywwgZQVE8lo++8sWSUn
+1v4ihxFXXKAeXfBXkyP+XNKwscq0H1lz9CsJcY4ZSqY3CEhpHRtctGi8+i+GpnH0ng6WoHIY2bK
IzM2Ohzt8+sku4uCHQ2vlLxiVga/f5foNHaKlxSX6UBt0vB9FIQ2uHSIFoMvDrYse/jUjtYoVYpJ
UiobPgvSUwrjg5V5KUl2XFWe/R9rZ/PKyIYGf5ISLojrWlJMJ22Zwv4MXTDrUmaH2ineBZT3SdyX
BMwn+xS94lr4dqtWry79vK8IkADGpdv4wg+fz1C0Mxz/zP21Mk1ir79zXJNbhAm6GfPaBmhnSWtw
+Ri+YS8NQEnXn3T9DU9fKGHC5QWNEcp650FLanadGs6NwLXVaLeHctqg6DjSe1Im3UPjEvAGRx99
sJdNIS1TIrv3G2Q9YD4JyGLMJH/HaekpMj29p2Rw0fm04sUpTN8EQqLPvQ//OeQ18R7DIXIqIdn7
TBF9Z7jhvV0xnJLPAn5FrBWQ3qkd9I2/KboHwExWN0L5xT+vAiWeAB2WUdeNhhNkgcbOmfF4U4ZS
SkM0l5NjX8F+4hPwU2AAi83brDXOTeYS/XFs8xjds+3DqZiCRTmyU3DzcnUYQNFvH88YBHR7XLse
JMxzeZjOGUuWGiyPAGwBHn0pX0whld/j4WHQGQdRo+R9iTagpGzPI7dl78av9hywlNj6W6uuVZfN
75E8tL89Riyw76IRNCsxddmGYWU1YpdC2n2ExKcOPiJM0x8D198jIc07HEvyvYAlA9Blq5RABDjb
fAanR8M2HUaAjUhIxQ+N7q4EF3d48ENVo2Ce2ygG393G9Pndho0YDmrIj7TBKflgHsUsNJNWdoXS
tx6GvQnwk25Kw6j8udJulahz2Eg2YU/8+4fCHsji/WIXyJrLW9sGRS0AhNZrsXHQyRmaGHOUr+ue
cY5ythcBAauV9XJJcQV3V87SrlXc13WlUyG8ntq9oB9XDItaEzJxEcGj1dHoiLfdOZOfoD8C+WIu
jRwAk4QMrv+mdeMijHCQMLpep5sCn1/cxdqn+bpsZtjbGFM/vCr3rSVqbs+9PZy6iH2kNAYOSfhe
9V0wxQ4282JJ3AbQfob+P/K75bx2fYX97YpF61u7rnSzl0z7BttbLpQj0TYJyNPVaq4Xq+W9Cmcq
1lw7ts2LhguK2gACSpu5D2taboY6WHoCQz910Kae7me95zirPaL2fyqGkA+h7qjmNiZxnlwAwdOg
W65tnSZiTiWYfTKFabyHcpRjmEV1qG6prJCRbhKi+a9nI2pVrvNGCTYFifyXAwLgiVuM+cdO89o2
fzS9jdr2XAbGjIZSZja++385MDRQnqgHpLvz7xtsYC4XEihxK4vefF7KEvZWl/dvgmh6g3IrDSjJ
xrAKe1QXG/qFJW4miKA2XWrPxqw6qNdqDsJ/dvPhRQNCbZC92L6TCCpRAQjYwGHRoCBnFiWcDGyD
ax4qdYugrVL+7Hg9uw+PSMbpBN8BWtw0Zav2wVxYnuDZDdjGvMn75SaH1y39e0avkYhXVKzRGzdQ
xl2Vxu4RYcf/bAb4ak7/pi7ZgDHkCmv/vRPA0YixTF6M5bumIn5hLCedV1s+H89fFcCDQnvLToHT
4vdjpSNRmCtt5aERlhSziwB029E1H5Gir3VY2CqkoK2nNXha6IIjzK06w9w9SXI/Os3niG/aRmT7
J143Aac2dq7wmTKDvDdOQteafy8BROdUEu5Hks3GZXneTPoEGy0yPqJ5hyKNYk4UZCPHw416279h
k1S/vbJZLv0hH5nXkBU5Z7n/91zE3Br0zN0XbqayT19WR0ygBumf7/jwI8s5Pm8cbzKIH7X5SLPK
E2fliJkF0RzUc5XU5iF2SoRN5llmaxWvOmByQvMxyQAxC2/jd8W/KVOvkvuCepoDIcLKuzbd29cI
oJJ4MeE2xk2qvD8faJRY9D3zBQ1niTXq9kPGVZzWZBmTp4GjPOazWj/mV+UBsvSB6Gp3FLPF7Oyd
Zr87PdbFqdMp6RmSq0slfoCybVJn7AUrSW+MRYjDNhR1WhCELiuQyDXQyeK/SqkZF6bOQErtgJrd
t+W5HQjjyzII/RV3XXXuBA7cEIIx0sFGTwblvJHxC069IKae5L3MlVu5CyPuhi5LFZ/vL3KcUu61
PYqbZmJ8NzZ91Hl62a8V3HGUcco8ei1khgHbPE7/08mqzCr9BHhd2OD6CE2kHfRe4BZDzwvXumPe
StcLCHX4pqLTRz0mYcOU1gxHGRIMEIW0aYx3G+0ELke+s4M9D7KoTI009cJd5rhNZ7CafelLFir5
AhQnszxOV1XgVBy+fggqRAYpeWqAAzAjnMVfOad2LJA/P1KYCFYY+Jhbp09+uOzkzsr21LJUTHbQ
Tj3Azg1CYWl/lUEyHtank0qLigfQ+o3UGFJSvY+YkCeiyw3IxGn/I+MGsKCYiDF6aiHUujkezhta
CwCFXokls+qc8ccDUIv7N/wi4nKNmNh0yitnFJsycxBx9WMMmHB3ZlEiBWGVJzcYYuXWcaHxvWBG
g5yE1UvDGGEfE8SITQ2OBogx7tsVB5XwYBKJiSVEDNn7mnlFLY3ynABZ9uQqwhLrkpjzyYHPvFsg
5Sl8VW6izuqsGBBg5VzUybtVhggH84cDqFQ1c344Y9LZB1v5e8h9lA+SpPNjhxdBe5J/azwQrQy/
6l8UqGx6OoBHnNMa3LEl8fhD2ODbIp1KnJ1ZNLGOV2P5hN4+tFSwMfcCd0QoZy36V3mEUMJW2Hxg
47A31MVvxGz7y0AL15McnyhdVtclrZ2U2gScDZtS/T7y58lGGvR2H7iF1csQ5E8zgaqcFURX9Q9m
zr5HL3+2mJSb4j2BCIeptePqTW61Kjs4k41h7MqDdBNofEHyeQY4BuLVq6AdndlK4Fji0/BNB+HK
8YBNUl2aakoptHpEbFhcUrtVppFiMPw6AyXGgnJnlDy6ZuEjIyQtYWRwllVuJMcvaHH3VzxdmLcn
5Mq+wrI70RsR1G5QnW/hxwHQe94h2yoH2tDh0u5/C2/5+ocZDk51WLZQ3CnaIi7aBZYJqbvBvXsT
KlPpFKuGEe7uMnGopNCtWaV5sgOtJPtduYwwVbhkxFVi9QSu5BkDjgL3Fnfu8MVm9D8D+33WOBfG
HCT+BitFdOikW50ZkWw8t3+CF1KezK65Rg9P4e1uTlJNkETRSrk3VcSUEGFHGHmroD2wz77+CkMb
vLzbuEdDCzllAnl4Rn2lrcc38dOmbWEaG4RbpqBKavhsz+7ni9SkD8CvDuN9BtXNPNmibm3xGj9v
SRdeXslJ5lWeSRi569IxaW/Nl96mWZ8CDXxpQmsQttemH6w5gL6dIljEy6vW9VSWVj65lCXwvYVt
ZCa9GXQ9Nll1GPF677i4sX304RLBrUjd3ivnMeFAxhgEO74IO/cKHKqjzJ2wXRuiY5lQBlcMlw6v
8zdUNNy1SJhaXTVLT+QEwwpz0PDQdadZHLBrN1HDMzOYlAMrI5oqJKf3sgfSxpJvXJxarRqhwFHY
ItBjkBWvbFCyRnog1pCdEpNadS6Zrhv+rqdNkv2TTNG1RBafk2NhMBaugOR9Qxa4giaFl+s+ssXp
99bIvlwlh17KGgnWKa2YeyDEbnOvIpDeYyD28beJRlPjDY8JJMBrZCkIv8ZuteFgr6orj72CK0fF
nB1YS+KrpDGoE+4Zhlyl+ZZrqEizUhhiaSTHdzqs3DV8gDT7davL17BhqgvT00ekWVaeV6AyT692
JeE1D2YYmAWitM0rxTce0Du6Mc1tggEutumKes9Sv254GTTLt2u8hYS2BsfNcJk7WzAYmzrMGdcC
rn2dUFqCZliuxj9Wgx9BKb17EpvZShDIWH1Mt3R7yMaHlTP8EmBr1/FsR7kuspeMv286fJzyalJF
qNGexVOU21Kc/PorqTjr2T1WDU5tDHOeJkN77avflH3+q6nA2GGuFC0BEPJmVEFzMFVyLI8g8zfz
0igWo7ZGOdJBRxzt08UJUz8IeAUMLI/sVAiCiy9ta+Q7yYizxrIbwoolBSdYixH0gTbS+1BFNfwu
xxTIrLBNXO887h5Fxv9bRXCKm2PVF99H0Ea545KdM/kKW7KqBhRRURBwjIoHfNUuPW60jv4KHbvO
H+qvAv+9Gu7BM5Uv+1ymcCCY4O6sVw03v/gFttygZ4pRhFMoe8d6I22rnle+WnRPvfwmF3UiuzBS
Rjk9EFAPNkbt7o2ycI/WpjmyLajrqPWy3qgNf0FDCOjzX6E5BD0cy1cQwZD/ivKi+aMVEhyQTPGd
SF9eeDKjXBTD3saEHe8KOprTkvToKBy5mumCJL3odHMAPaUEk/vQepGz+qozqUX119Qy0E90+U0h
7/8X5wWG2c8M3WYDFtDjNx93y7L4ZCuMSMLB5HbdHI1SKotDwrlXdkcnNkQToiitqez4M4aSWoYE
Zn85fANc0aKYq+XU8eR28TryciCzYhzuRrpAvqzf4J0MuXFwhUIXfcc+vEAt8nG7JSSHweLnJeKY
x2F7IfUELATAQsss+oBkawnisi9zy0Gd4izeUv2gFrSVy26ey1f3oH3W3uG6mSonir2vYm6gV2Bh
3OF05lZSQKWdimKMXTfkVaXDJdbBOESpRlDLAVfnuNzs1T+mVFJH/ETgb8MZH7EE7A8nr+qxsSrq
ULMUZs7VsIa11u+t16y3LcKGR1E9OzQvPyMYe7UWVrUQZYCNPhbMaZvE1/xX8sOrtHq+0iv+HAtu
LsCLYOI7Rse3ZlaCucYbiuN3dFAmzbcjedm6BZPOSCLD9e+AC52B7ii7FRGKU47Vej+/lAMMsBrn
1aic9V4wMW/6CBP7ypN4rfl7OPQo3anOC5s0qrmHoiEiOaSeiC8uXPBXzZtx9URny52WZs4DrxrH
m1wD/sHPEuJi74AhZwcMK+wBKwpemeUgDhJVdzDI7zQqFazhh4ErMXWd+fkMur9YCt2n/sOSiQWX
FAcj+Aisdou9qPt/buSO4D42eX3KpMEsH6/OKxNiwIvN2FnbGEiIWPwN7DU7u5l75HP92ZFdF5kx
t8uGRIwdWTVRLvPMy/bxRjICqXf6YusVzst18bUIEllUFGRSzOyc9ebYrC08qHVdZBH6tyOgXFep
I2Sk4vI+ziX/x5H9pBuOyH5ewMYadMFifxO3YDp1qq0DZXjUwuFR+v31e9uMkYY9aDd+Ip5wpljT
+y8GjsH9XVGsugzgmeMac238V51aUU7urlfzCo9LScJylN2CbKW5FDkSi4duRQG9VTbHjaQwEU9H
XsysfKuO6+/pO3oX1wss0HpYJW+W0ZNKtCEBMLimacqyZoJOBdDphH4rkTux5N8LNNH5oMcL3vDk
Aoz9L7OjvfAT9N0Zsn++SaZ92/hCRgwcyOWTIllStMtGycFX0Iqi9iMGoFvVjGNUQt57bKT9bSwl
6DNw/uC0KE4EBTJWgYygCFvISKEeSok5Zl7yBMGL3B6BWS9Zc2M7ewqvnk73dhvIKvkbM8/ALKQq
hifJUeNy6/7KTAYsm0CH58zkEPPzAIHuppZJzmgkpa4uDSr2XxjnmpY2akADIBsz8Z9KAvoRrefs
xlTDEo9WsbFj3GiBd3cKhFBYbXTUtWr1l0+8+pdXdXML1sjwqij5tY3K2ejIxk0+UYSUyv+v1z88
02aXamb0xdSsRjC7qoNtVqBgBYul63Ud2/MQce053+JWkcrwu6Le33Ezy3XnA0K+Kv3B+mhtAsJ8
RKAWQGGf6PN8nQTMbbRuNijC+YXGsLm/vzUil+WsTfTFe+pgPsLW7E2lwTOgv40bioE+oGDAtq8s
+hsZu5X0vJC6TTVnvOCp/o14VTCni1qHI/L834PTBjbNs6mVZdhXVN3TVdivoHYCPrjpyB5kBPH1
jt/7+faVizQnC0fRw4whUCdEmhV+e9xkxq3SjbQr8SJVm/M0axezjTtqLtWx4WasTk0nvb9QRthY
JpjSJT4LV2uoSsGvY3NtH2oXeC5W3ZLnOwX2/skst2NxY9zoE0H/7TwCsuOpLbEirAsckq4/JnD/
el9QmuLVhVI9IKSfzRjX5dqsHaLWcWKU3DgsEUxFWV86fDprflrhQ6oV4dJKurlAlXJGMv7CQhaq
zMLMxK4MQd+hE9cSyQVA4V6RM2sqFlxAT16XcISD4lftq0fBygV5AzzV/790l1FpuZ3PE1DGVL1t
+y9Q9OFKaKZ3MciuvN5zOCpygqoDztvKRmdC7Zx3cVZi1MrqL7nClbn92w3yHC3egUa9/p2YQz5g
rKXVwlp/xY2EBtwxNZeO2kizU3+4cJ/HbO5vWZIdFoELZXk1RA+Xqq65wSaSXgLIH6WmHi4abcIw
HTTszm4NeiTIIeQOOpaZpYhXj5r4P9d3kCzTxhsGQwztl+KjUAzfB2H42WDnTfNbJ5aLAnHUzrqK
38EAQ1LmpQrw57U4COOKEHI2ka0cyq1XogU1CMG18IEVv95ozoOqrN0N8e5m+n5nPIuUIzNzGzSV
4SwLEx6Eidpz7mp53W7eldgTbWWnwfVYgfixYDoKt03FoI4EE5PlzoNiy5otmt4L3K9Wk+z44bWE
GIE0vH3LRlgLkMfOaSQaYgqgtYeFa+WlX1gVpkxJmo+XUKzcCB3XM0Qj14/BIDUbIXh0YndZBhjT
MOBHFPTme1XaTiseDqsIg4CY+FGbxBIkg1NiWqo3hsp0T4N4XNzNMctUpo77xg1ooQ4jdVHDkJxI
D2IDdQih1ew9k23NAMWZArlMqDVqaGNQHjHI1ZOy+/7z7LuGNWsQpH+r5eDTXElqH4HHP08Pre18
i27rJxnMDVlUEn9TxLAdOCbr3xBPMJIx6CWEYIywE/13ONjenlTnAxqJkahUMuOmqpyxZ7XmzXwW
UFPymRCUXJh4M2WWxG0GiaXowhnnBXOW5AP/7LW1RNpOstT0tc9RZ8fRj21jv6CL/qPSI6VerVTP
BzwH0r/n8fMF9mhBwrzQL6nwe+048W0uHYTLP2devkhXtz8Py+AnihovXOBDmw2yiebuHTBlhLZY
0glGCyqF7Cl8V5eacHgbk1aDiXSJ0TDZ6XTd40xkh8O5yHukJg5GUlJZh4o4jCH/XzUtu49/2TAW
ZT6QAU8ibi2z3TadvMZZC74OjHETK9qOtCFdCQVDu21aOuYd+nAwgGEQhvG4l693RA7mrjtU2SUP
RDJMRSAy4zLQMZ3TJfOA2SNkf0ldsERWTdIj4Ad0RSHZ2MAT5UXElwc5VeanUwlMwQOUJHML57r0
w9QDPOOWWpAS4RvBegTZTp/BrepdMIIMyt7glx7CLJ8nzCTDPiYO8isC4shaGgXZVqCopDzaBpFT
n2viH2bEVyzlRUeCeg5ghyWq8ZQwwaRrkNcVtPjYRvBk0yiwICI0Wtdh938EZrHSFiEijIA30ZMZ
mLVzCUytwXERWdOkfokDT9AIScoAkh5gOhLBbg/BOcIuSl9P/riE+SoejsfdueGD9X+czPobohS6
O5MuToWejeETWEYlV6QFkSOOJZL4/tSgVQ+i40brvoYuGSK0FTbrrsmGxP4oSC3VtxHa3cqI4ZEB
+W+UpMFDUtO3boUbreVAq6c91LFIAxW0zNaY/nGVzxcZdpuY/4e0akJ4pWShv79p77syp+u0N2dL
Qs9SyY3TJlOqzMAwJ8Ir1yKuCEbeLPeyGrf9AhGKH0nCbu/z/MuCwF75FFSMUNGHfE4w9C0lDEwh
jHYkA5G789mbhO9PoKzjrzxT8IYK6cNUkHB8bSP6W2dhC52kRLCmCdUqC3ZMJ9IO2QzwBWVCyuHU
Uz3tLc3gWF6Iexq6g+otFns6AP3S3hbP8YOZvjbXTi5XgBZlNvLGrcMuQORKQl31jKX49mRHOYTI
Wk33cqdXFHX3jJ9iURHytlp3xQevnP5P9rPUuPrbjfTu6YBMo4neqbphHAFCskB7VNGGaO0RNYBo
TRL5QJnV7mlm8+dvgyTHp0saIUaAp0bH8dIGwBUQ9NDQ7PpAOtlI+Ib5jOalAcIz0k/NENcr2o90
RKIWpBaN7JpwQGa+kHOltLhlNi39A/ET5+rN19Hw4DgITTA7s48y3rVnvHAthCC7JtMHCjHTQqB6
CqEu2T8VkElEO19cvyIlqwIXLQo5zXBm1+lbN85z4DECLYPFlY8AAa3eXfJKFQSkUcgmSpzLIC0f
ODNtOq9MebCNgsKlAcOiESNTgIoYwCUemID/WRe0T7bzrcm9duniMtArupQ4AQMPbzxJ0uG/N0JG
iPsIHgN8AUvN23rYtfxsQKRiu+K8c1UsrhjRPkwMKQQxle7eM/Tyvq+ABNIabrxO9+22clqxZxH+
D1SHIWz2YbgzvpvTMpuaOG/0P9ZrK4EFT/6WiZpznAuClvA4BXgH1z+Yw7+H0w4eVhAiQFebmdl5
C08aZcABawfmcq0eijuaXVf4rbt02xHe6Bay4J7Uz3HdfpghYWSVgVIr/coYBuIdesUBuOqhiyVm
uAsSGaEcEMawOQk+t4MhfyID+Ni656odNjdLnUTGVNqSgdq7rFpmtWQPuozLD4eNy9qVHTTrXBa4
cLIXyeIIW7LaJ6BAyRXiOckxYFFximGQ73YHWev8AQ1NM7+wfbA2d/tkSB6c4msd/f9oWnl8pyQb
Em4ecaie5lRrS5TzazTWQ3quNnuyJjqA0qYjRGVXhBif19KEra66eBTSqD4HhrSQ6jdye8rf3xfd
1SBSS5AMRFdZlwmaJ6psIOD59C4ovbMGNQJ6II92WqPX7+2WboWY0NhkV2FaKpxwZWWbkaJ+FG4C
WwCqCnpuFgPGUxRqMp1t9moliEEXJTEJQhZnot2xXYO/Q1DkoW0oNaJloWQD7JbaLYix3g7lk77x
j5tCD+TNb9ZKgTHSFurKuEMpV0CcLQagG7+YkxvXyymBtcq0y92Tm0gP4XdoITARQ2GcMaay4gZ4
VmtDv2mXgvZautFk3xOwdvIAhDhgatXyhBsgZrIo4+01ppAqBGxFjZFJMviVqGglgVuOg2n3peWf
pUsacsCKimHqZScMSiypMaaidAPSsddxS9hDXWkDBYstMSgGzRncYR74t+RoHxIRZbJ7tSpn6LAl
s5ngTdT5EuY+UlJPR+vaoiiWJZYcbChDJRnu99UfNo26FI2aN0u20B6Zn+gDWSHvnemyF/4qgH5B
FCkWmzIGc+iicmdL29jKmfQvsVm/dJm03a42ElsGn6zIGdGGQxH0FDKHoUbUKGgLvl+Rqhm56LPG
JqmqpzDtpBmnCS2Pffw9kxy+4a+UC8RaNmsAAYEXvezxtHoZ3BvJ9Z934+PMaxCkV5sK5XCZ5pKr
otxTD4fCbAmRwO+gCSepC7Jwj1VNs6vot1ags1egE8Aq7Xc+Y4krOir45/Nf2FNXjULqkf3T69oi
EH4P3HIxrsiZFSTrwbrlbXELT3E8SWJ+wWpGnfbTxv3m33bPAKl1arsrKSUu6pD/VCQkgSnZkxc1
9RcvIedifQ59KZyc6c281S0KTWf2O1TWP97HhMspoH3t8RLcvQrwGC85QvV+iMlS8rKMfLK7AQTn
OVpCZoaexkU09eJ1CYbukr90u6KM3w2NaLsfnTrv05f9ZSQ6WYfsG6Ry+IvhWXiuba3McA+Ar2V/
cqcsFRB/reQYJS6B1l13s1hC5NGWqHEJAyVynH0y1G6VUdosGnCZpmMZhBJ62B7kG4IfLpP1ojCV
5QCVh3giqNX/2yjjoJGfvoYW13myqZCB3PFzPDDQ1hR5RPEu2b3KxeqTg1eR7Bw6GDt2Pz0afGOj
6Ob3Q+xh3qMhsXqYrjfyjkFeUyb9rJQj5BRrwnZmktWltBnNoNiCDP0wwaoGfWu+w41U+Brmnw9f
AAP0i70v9OtpNdXUbLAXQCi1NQfN5z5gzSq2Rg692JOx56lBFrzwAOOykcHqxpmw9M1oJVUq9SNd
220grP4o5dv1bnAQ0+Cgz+DyuYwEnUangSBmCvU3EolBgSPecYJW9teUba7j9AEpY4LFTWqNogmc
70PgEXxr+jcBxdJh/pu+Om7cXsLtayPvo0bP9vCU3O0VuwgSHfos1KmPUzhyFON+VmY+Ls0flG9p
OEZT6YXprkk3UOLMQsT8CNZnehZGpODAzvbzH2augwI0Ryq6RzLXfJb9apHd3N1lDyLYHtF8noW9
42myaV07DEZQQZf5PdcCr168P2vkArZ/np5MjGbui7Zj58ToNvmn1MHz8Je2IT2pE5xfdvpiNNpT
h8eBhOOo6WdP24RLgCWWhkYXvuxL/+I93dPIT1JeNMtq9mlxN0NGJgLmVkg0ZjEf/EMP1nJLzMrw
PSx062/R40spIxp/0bWPUhSWpGNBCUUeYZkQ7vZNRS4KXKLivgoM5sxV1zE7GTreRU6VZULU5eEc
1Ph6tD+wAe4tJhCazNEJKU6qFqJKUcyBgtEyYTPYhtYXB7vNPA6SFOUDgkR2sVSqYP1gt91KhxQj
M5FW6Xl7Ll253VtzHeeBKym6PKNWCZvTXGzFOqidEN/BxF8ZbfxXZwssJjOQk25XC1ZDQxmvVucW
UChA9pW8yfQ3YtCINcS1FjZP727pa0NfJNUKoaJg+9IvBSFLhAUraXPI67Ghpf3MyeAqjIeInk6C
8tMqD3cWUBtnu2fO8WuQ82KhrFAItCQTMFOfX4DjbwkJDsOjncIWCbSkmN1Xy0MPUwACgWC7lKLC
uy83BSUtS25GjW9FJHsE5sa8I6ASWBR4oVNXegj1VHwz8CbicFDtNFu4pSo70B+YK3n4GnLusJVR
H+5yOOKo3WZVHt4rMtW/lV/q41uqGpPyObBufnuiMsYb7auxEHNfFhETyNp4nUSzu2keLYS0azi7
tkU79ghl755lVDTzE5SmX5PBnaTQsKOX6v/TAbONdpUhfD3saB4rLzjVuv7kJrJC4mt9lklyZMYw
J1jYMtxyW3atDn9sUggztewyZufjg+H7ccnwNVbWT322gZ0kMOJRa7YjqU4Y8X9NpGxfM5FpyIag
R8lVxsEG+ILkayMemuM8+RGRtt8jEDlN9lRyJjLsOmc1RXNFqzZ2uds2EnoMMPyzOCyMB8sn405Z
YPtO09nSPUfSadOGGKkNy6vChlNgkk1a3Fx52uLWEzY/UfE3T2Y1Jntq6YYf8gcN4MBx6nZ6VELn
ie4dvmN3z9Oe22KmOCUe4Is7i4+4mO/adFaIciOcihIFJydmjpIaRnZeGTSINQQ7HxffnCxUJEmP
1U3CwZMxknKrghp1yH+HX2YMAKJNUuoBEISSWj3f21a+7KjlfcHSi9TVk91coR731iKapnBwGgnM
72dTTVN3/xp5RALNqsLxi+CywbDka/2MY2O27i4ob4MV2PyBspNrbItJIzZRubsTagtk2yXmvuZj
pdFTnvbcV0X4lE5tcgXQRGioNmZllOu1D/SZ8Xm3vRQvp2bQSRID0mGxvHHdNAJdyg3dVG3tTvX8
+zGVC/FOOYNNa6Cck9ZJInVsmUl7JPbhTKvr5N7JsCZgs2d5UfAeNNQpW5PyaL2Rw+jZDoVXJndR
JNfqF5Tw+5fvw75wwk10IHU2tUu7cU/O51Ef8ycAGnyUIEyiSVRStdcvqduKnJQin0NAHIRpXnM2
wD5tm3MgaCfcg5USgDanHduwt+mg936yofTSHo20Zyeol0QyNkBVvQ/ezFsoumaTM/aubUvfNykH
6MdoeS5z0ap5j/paD0pQPof4PCo3PmsNTxVBhZaycxgz4ghE9zdH/FFwY6VU0ErU9VWll/kkjtdr
NyIa+i8LvrQLzAkgP4T4htZA+h1qRjea94wqAOX6sAD4vgB4xM1riBhSxRN6ZNyh9ueUJNHUPdAu
AfYLPhKPG4IJgd1con3Jm7FXp/eI+yb4XGO/FBG/0OmaVBp5kjcU6ipgXOn/iGdnyNr2tGvJBKVM
/x47hePjQPnpVPa71NjXyr5El+Bw7V1AabT2Zz/10qqxYKhlHUks0XR4tquiDqG7ST6dyd3DS6Bd
xaJvtAcvDONAd1QO29JJiOR0SkFLmKn/GJ2j0srpnHSITmURWoqfVZk+o9jtzz1JFYVrsDAKs+0B
qY6wEDYPwsQyvHktGzZM/fxviEt95ShjlqijvnSr3EblKFrheWqLh/G88r0vs210DnNrrYQeze98
bvu298pD6tp9fyRk4dQK2vjPclhV4/PwVghg6Wi+2RQWwye4mMOL5MKV0r/87wwOjQFuypIAKzSK
0rHwvUjD/NGaiYdZ4KmK0XaMg1qgbOAcTbmfoP2CptStWY8LPAPDEGbdYtGTpKltFzQ6ltzSPOIP
HDsict/18D7OsdWI37T6PeejuF/vqWjq6WBnj4o8hQ4+USSAd6I8A5bOQZ3ehlxCnHaMDe2pr3MV
IbbyGPDz9KOfdjBjctv0Gkz16ixt7T/2qWMIeb6A6XE021mhQKnjD6rEbzIYHi+hm82P4OiLNwps
B6y6B1Sg0J+x1GYhWmsuQh37I9e28joR9F2ExJ7qgCsyMEs6P4Xb2lX7z0ov9QSbjvy8mInr5fTS
YkipDOzuodBv439nfZ07WCuGDAjtUdltNLCTr5OYOADSt02Sds73hojWiV3FfsMB5Gdvs0O3kIhV
0c9rrEChvtzQMVaDjxo0IbT29mBnI9f5yPhpTei1EJ3Gi4Km1nCUS+VAkQS5Wi8v97oWe9WfWeVS
jwN5JnKIu1WAtZZIkUDx1DDC4lsxFtey0g+6l0V5M7neZHxf3Z09JYZsa6VfY7L09yT/w3dv9x3E
qWo4T9IG35XkqUrcj6ZkZGyCdDBpJ3Rx2Y8U6bf0oWdp7na0dqEqsy2UgB/WuVARzakfCmT3EZS6
eGiZsYrNyDGEzSbSin48xhxBoJkqA+CQ+WLKd6/Td0yusC/9JKUFGB8tLGf6wTRIWLpvDkwqRa/d
GxxxncRKnscCw3DOTsTVXkyI+pWakLg76cewUJ2htrhgBm1bJZpUnmc5YDkn6NjjbQtvMYZshfV4
1d0i9MKRyIOBykYjQF1XodenOfaUEJX7ZOvmmRGsPhFerwuWt4HtGdMPOtkrPudJG8mIaEHn6urE
WEDivpfuOVCHUC7BqL5jeIGPhQz6MGCijpUMPaEC+B1T5VzOkklFssMH99Xf/kYWdL2bwj6y27n7
X4ixuuyDpRfj+HsvycljRwR1+l9anp6b2jHlMk9sAyhX2ogguE9gUy9sOZVDpaHcc15xfwnWHgyh
0lLdWEKZIo0+WuywfKnr51RhFbr5igblmvVk2Gw9OFEYAkmhvCVYSvNtYbSavBRlWoL4PEHpWsFY
D6LpfIy+awJx3YwLCX3tN7UrrgJ8l1A+RLZZsbrlywaWDhMN87X5KZqLEdQdVhhWgCGonYaZhWjw
ShcEAzYAmypUOzHy3V9TjyuHPWNgN4r8UZiyM/K7dFzR351wd/OHdzbzgM31GtN9TOm1Qzo424XC
SPoTVmHrnDgbuV9biZwNkrRTKbOV37PriPeu054Bgd/PCB03Dz4gNPjINd47qsEZ1fcoQrB0iugZ
MW0odW1soQ/xS7Xq8DlyJY+2dmgfgKhqp2pQmVp2P7pFWkdq/7HgJmFNkdzmpfCDDM8Xkic1EQgu
ZrODDLvX1AVYdkDSbScprNA24d2kvOsBp4oQIA+qIAnp0wd1QPamgHLlft3TN2XyL4Q7ZWjxAL4s
qbFikPqRtENFC9G2HWI2e2Y+Nsq+mg/9dNwNFsekybCeqvXzH8YNgnlJ6QZTv4NSWeqtKeKrbm3c
GbmLkH8OvHle98WMiqDZWXNpLlkwPmjp0E8Qih1OygyQP+Dfk2ZvQHxXUoGM5aEA1chBFbJfFbD0
KUlfDhphwmUhV8iDLTJEyj5r9JE2CXlAWFr3c4O8q55F/JabmGt21cOS2UdEB1LOZ6vfX1fMil8N
VUC7g5DRFnn8nlM96aWByxn1d7j6TUo4T1Nx6uKUEbc48Bx47uTgcTvxuJlnkhg901qGLOH3RRmU
3O0Pw4gtseEfSrZGL4HVrB4Ertweo9jRM9xOzr6As5dW2WNFimA/Ur5zIByu2Z3uphnQupSOnY4H
rwTMTe5HaCFDFtdKCpfyUk790VjOXRvvifsHMsCL+JcuqdX/CWo+dHk2RofChJ8QxNGZ6GEQWc7U
XD7JksMQmT1F1q3gS4h4SduaijkN9TsvXSDzcZnBnW38yAhSsN7vi866L28nY6PwlWmhFFWQz9Fi
EnzNWx9pJnJ5jcCZ7ggDh+50SL+wJcmLCraAh1gPFUje7a2eKnA+FoFfW20ge/yAOB1CQJ1YCX67
HJM/v/o5fmSJHhpiBLnCBfJag6Q29e8ho6Ax+urekrQhsKpXh3/KC5LzXScD2lZRk6QrluCF9uN5
NFaB0JsvHG3viRIIcwl9lEI4Sq0/52y7YqKVcECzYWAZYo0+HGpGnmAGDkmc6E/2LnGNGEKoEm0v
iM6KbkQpitfb3nj8XUYk0mOSikBDOOgc3P4qPfTZzUr59dzExv6crjzvmsDptU6gK0Hx9T1Smny1
fgcDBL2Ba7zrxVW1wzkUwPCI7+pDlNiTGsRwwF8xfVLew3NRPoayQHm32glucq4yUXdN5wMLTRih
iZKObivZ9kwGfMGf3GwYu/wrTZwJrDeVQ6+giygPHwpIHbFqOMe7IJabdj67xiNSz2NLYSyb/Q0v
VMj2NMzO2FlpxXD+SPdyxMbiisj3AWuIB0vCvOL5XzawZcoDkoJ8hvuPKhmFmlcxrm7o2eMa6UNt
V49tU6Wgs11mBojJmso5QklxuO4MuLfJbXAxd1hNYXLCUJEE8JydExp8NCmmnd61S0YVV0o9Q1aE
Qy7KN8on0jK1bP2EJOoc5ns+fP9kqgTGVtbGlBBDu/gHOvX3Z3C0EOrNyG+8kQPUxI5ZdJ2GQ3lM
Y+D4Tsw3FZnTw2jMmWF9mz6nKoeADetOt3CJMD1Ng1MXueKgFu/E6ZyhR0HXI++m3yvyhj8ddrGC
2jW0A+YP7K9D7ir6TxkjCzI0nzTw8VjRAMmYUEi31Zx0Sq2YlSgh2hMaixV+oaNXpiMFoZHll+bv
/8kjjwPkoUAven44XWFb5Dw1CAhKGXA0HA96G4sHi+4BqEo0kEVyhB7wb0e+YtZkoKIB0wabMcri
trjRaHdIcqig49hqAI1Rhw1njnnYyp6phPlE+h63vbr5X87PuFoN/VXfLfVqCxkUR3hz7r0++MZz
Z7EyjbQPkj4WzFTXDH4/daOZXJSRkJSpDJq81+JQXvrhcot4g6w/RW1KneEBrfpSGSDvuDnZGN+x
+U/Fcyrm6/DJHXHCg5oFnyJAIfPZUPKYhrFTLbzq+lwnRh8Pf7gvXXkNlEQ77nBzsTjpWrRo2Bjl
1gOOgKLj6DPHzR9ADQfv3DVZGxJRxThTtwTDx+Z8F4CWtEauiUeyX2TUV5x/MHDr3CdRF4AK9glv
9XZfRh0Bpx7fOM1y7KUBR6SVgJOaB7mb28FejX2eHPfbfCwq9wImMKyEpIqMUQqjueToCopI6ZS5
9hK/VcrAsvDMm1PYJLN9Did73Z9wPOKb2g7NOK5YnZCl7rG7uaXmETB0Lh8/glmbifAL4TeeXZPc
2KDZafZOC1DPfAwlf8TogfbZm09CrhwxpX44njvEDQHp7ccALqobfodmLLmbgFqq330K5xNpFycA
W4Ag249NO8M6lr7hDHIvol0roLQ8Xu5GVDef0EK0As/R6q6lsGGoQ4ZLvcFw/Tm3lLcmaswI6rxm
8VVcvNHwiYu6rV+1kMB1Vr/vbOlH+4+iu3Dq2DeTGLuHwzDyNKl026vFCLPMuHtSvi8fZ8Xb5JyV
FgnDaJe9gnruB6lBx2TZYYEXy+gRTGZkeDtEgAnOEpB1Nama1f89wTSVsHSYU91dIgtHDtXx4bIG
aB5g1Io3PmLmEIuu5lhG2h7xorlamssdDV+dgp8CADfPNRPfRPyDVhg21vCNbAQmv5e0NgC8oSgl
FNaFeja+BM13D031NT/kzZM5jjQ09C/hyrGDGNc3wCnV7xiU8+xX6mVHR9ei4XY1rUT7lf4LAZ5Z
/BOKFMuuKzJBPDwMra5QjTnu+LrjuRQF/ajqXmqffovDkmDh3yaVaeE+vnudRWCpo7D9uSGSzvvq
Wzs9t/c2IxB/xnIVGG09Drb2yKzd/8f0Y3DmH4Z+fgflAFDqZYXNpu/w+ZeDYye6hc51RGJxCDcK
zuVUeLm4RqCxyGj/RofSwKMV6ex2jx5gQl4Fs54w/vagfXEjeB+FJGsYfrprQm1it0oFbK7hYbB4
3lYSMhdYwONRVShxsZ3U/ZijlhsrHvk11pNT4irGfj+ig9hzrLhaY4MbuLK8kYWuimUSbtbRhCrD
5gme52AYYfrODrwyrYB2YD7Vg8J0Y00tOaE8YGwP270UlzLNGr4IbbX1zthtbPvmJvyDBbQV7Idn
aIisKM7buj28nc1mmBWfwZ4PWJVa4EG2CzwhcVUDlAGSpPQSzpB1VoHiKtl8htayEv+vwImN8WC+
o/cdDzKMRd1StKM29NDAMI/sifAImu/w6K7zUwy6tabBHOcd//XsC+lca/lBQllJGHbVrmoGGaDG
9NZ2/hmERLvJaaFj3xTM8JPaMtHr4T+ADodX+35hFARQR3XT1JbJotuCtsqMfI3bdF8nHK8gzcNK
rl+HEBdF2uJOFx+RGiajSatWScTpkuJz1WEWCUezY6LbbPvUShAsxB0nfJ9irUhEytpHjrV8d7yZ
UAfebZjgpdzKP4iY3YMCgEV3PTw6/aXDObjbl/iyN3h29f69L+yqGJ+At8fCOQq/PHYihviZ9GfL
RFubDQ8Nxd38cMchS1aBUzrY7IyqI8l0t3KaMMQTVqrX80jRbqTDZhcHfcQZ4eA8Q21x/XbzUO/Z
NYpDbHZ3vEy6EjrlvRnBvtnPScMA2ZzOLKi5IxmPax/1esEWw+I+nXuOCAfTQDV0mzWeUuZpFc8R
RzMId2fx5qwHush+JkluRpRw8g0D56oc4RBF832Tb8+AubC9WbHeuvxBYFzla8sT4eQ2U39yDiiW
P1sU+f6KMKy0u9WLlNJ7668G8z4kPMkSdXKNRUlnDr/ecRuaGLHnHY0/Zt64wOjYXNf9/0sKtLkg
MPgaFtfs0bL8GHg1iCyM0awAB74Arh9LF+HQezHZfZd2VvqwFGzVkQm+otawzZAZMAEnwFRRuX/h
kY0KIG0GoXQ6AtBGlvpjARaa16TZcTlH6+VuAFEGpWKE/tutb8JCllngsmhxAlDmQH0NhL+6/hvN
eDD2PXIL2LdHCLbs+xLigx/HeCCmZ/vBcnIvtgQxR8ThE7N67rfY77RR7yp1EXF4i9h4T5e3h53F
7b8Wpjv1d4VvqHfeOMBQJEvr7LTlECZ5INO9+kPvA5iQ53p/KKsIgYpobLRNB4OMjtMLwNhdwIr1
hjbbJGFoBF0KyFYbblOuy+9xhpgrLT4Am3Lgm7k5T1nZHCA7eNLZPzh8KvqeMjs32rsRMJ1uPmYR
gShiE9xx6eilEjJpNIsR8Xqtur7toCN1Dox+C77FVr2WV3lYIMD+R6xZc41cFlQthedBdYfC53t1
wGQO3KkYALE9WyQcy4NVZSg/vLuBDYttfX3LE2o2I9woV1Fuol2mXdfUYQaWytFQeCBHVB1PsvIT
BSg9PCwyPEMmF/gWbvyNdYzKdLG5yq8ypT4fYy44qNm2T3vUgkehIlVvejeqe68e4LfRTJpaIiI7
ynPQ4MIDYjnDNHCsGGu7gLheW5U5EXtxkdQVQangRVXmgrrr4py1mXzbIDIpP67uu7WEWi+bDwGY
j4bMOC941BessMz+DD36h1imzzn0r5odhdAyeKuW/OAscP2Yc6zanU3u+qnV0MwDW+bPRx3XjaUO
hT8q92zRhsRxOQ3N/msyRp4NiPCSixeCXJrWdYOLAoSQAKjNorI8S8y2n8k9nhURVlEADxCjdZTp
oSbCG0/GHboubpM5Zn9Lac20huO1SRCmRzxN8YsUH0hDbup3JXgbQ5tqgt0RkNJy1IGGZBJmjtVx
J4JXzWcMMeSBaRB253PKmkZOwfZAKSmhUT9PnvyN1kzx2rPzV7EWXh6sTod34eGK9y4JbXyLmn+8
+gPNOrZilvQhlzqD3tEWXksiHMxrQ2esFfSjsCYC6uZRn6k1dd/C6E9Ybl+5PVHqFN01Lmxr0HJ+
U8/L7ijnARI2JESYW2ZvRupCXOxR5qgmCRPTgkQP2cvuR84HwwcXmVUDloXB8S4EDD8C3wNOkn57
r5jxWvIX5HkqIa3KwkY/2+eXoO7mGO01voZlIrKSgPBX/Q/gIOm+bpaBrdIrEG1Nf8CzZV5pKAV5
4xV72Z+uMOsDzP0nVNGJkx7rUR4dBuQHVYtfRCMxAjW8xnii5gbhMotElHxEuzUQUHwkVlOEJgl0
mXkj0oeOjIc4l/9oCcjAamKTL9tMk47rANhxYS1Nv8kvjCukLT6Et/f98sO3vNlY7YqxGs5NBd/e
C8+Dk6QAOWvE2TBD0eJnN0U1/hpM5rIsPqVuxI8TglRUtms60f1nlKmBF9qRvBvLTOyGm5FZGpA6
8AqSbTXxyZUT9Q5jAc1ltzS4LnbaDiXN+Ztrw91hMFX9iG/0qQGCJEETNk3UxGu5jdG46EbgFnfh
bH+o86XCHxQZKq16V/+GdbngS6d0hDmUyogMGoFnwKmo2cN+3BWF14QTSQdMVLAkJmOizaw+S5Tt
xGxYLxRJdfOs/kAq4iKiMFKEQyH933vvo4zo4ViY5nzBYQDeJdoWJVNv1UbF/5JLTA/Wd/9ICB3J
iue8Nl97pYHMk3AdgRKr7UVvdDwHTDtxJVHZaOw4WBubwCL31SXq1oilFzu95p6k13jWmW7pbZPX
tcEbk+jYz65FlFSGYsf3EpfQgBNrGx0FwrugxNWRr7Am8LLTVr09ejrR8klzn70uaIuqW+T5hVFa
fjGy+pIFiJuYSS1bIC104hAko+ODqJpHSNFSqq7zZvX3WNSY5l/PkraeEAeosubKo28V6qN2yIke
fC+wAUlGrcoDhwdLDNnk7cg55oaIj6a37GeaV5yNKc2SNLYytLi1TawSgQCR3gPrSp+dr4dQjN5F
rC9qJ71tPsqwxE0ck+21aG7ZxgjSzn+FzE4DvmYBEBU975mIt43+QUCaPlLVeLdH4V6LjHDgJIF+
Z3TFFcQNb3bahSlu/0C83+TxIF9RQvUbbbIWN5hRi6lzvAfs8Bc6oTj8jOrn6YwWL9knQJVi6vZt
Njl0+2B8IPiNC12+k6mt1WddtIyDigAB0oEMTXmbjPiB60bLs47zvhd1cjS2UsiajQQOVdNWYhyS
57DBFvL3Ty8fC9BmLWa8Lhzo8CckUl4VHh8paxhGCRTqhVoD6Ebe/kDTi24Kl1a/+K0ifcysx3io
wFPNs9EEoXbhB5GwmmOAAnltp2mlZWqzz03IMiIr/4TQsF4gpcoJchcoEL6iulonw2eONSAmEzs2
psx6RGh//Zw4jS0EuYq6ZxHHc+Xi/tG3UPl8fDjgwPAN4NpkaHxKS82vpOhHfaMRQSzLCXV7v8m1
mWfnq4oNaeCJI1YJYhobfZ9NGwINf6znagEqlII9JKu5mqv6/L0HugMcPCyhBLzTmAv9np8AQtPB
9q+iv4PNjrF9cV2iZXYls0M87T1fwKj2oiDf78hZdCJQnphojmVm1n6QVu1JCqTlBA8I0MoQI9mM
mWStq0SLuV1jS6/Kkf3Ex2C8yiZr/zgf4+RZJsWh3LSp4hIOEfFE5yI1V84irZYST2bZWpMFfOzK
m1E6fJYHw9fQ3N7KfOI5xRH5W5nXGL7pGwWYgfcSWONP7CiWSYtI7h86OLRLZADc0dpEWUN9cx8K
LzrjVqv0oNQok2rq2V2WjzKJYjHI8O7aKnuT3fSfksu251Zd72+Zc13eaWCDQYcBEmof9gh9Ai+Q
PJwDFxDbsSklLvXz1boVH9yJ7L9vKCsO35KXqDl4KhYZT+W71YBHXZzdB+FOzGpC6olLO1JI0xaY
NWpmP6uKs05P34bLV0kbXnKt/E4pr1OfMBaGc14fO6kIaP4ELPTCmX9f1pf56JSo4l+tBasWj7yB
5oE/UqzAgJX66H/ID+a+TOFYqy+3+yL6O6JxZ2uke47gL+QD9wuRGdNSC+nsxQWMOwrXkiufSs4X
Bgr/SBpervo4PbKjlELa8ArqkE3LZRxyoZQuGCRiARuudQBSHVbs265HJ73DmTcAghLkQ7PbaGuE
z0wdHdEE6Va3d4iDEsDMzMqG4FFcSq0plZB3V9MXqmGuOi+bLBhm3tXoSvspcOJ1hPiTg81QoquH
tyoNvLEKhqflC4tkE50AlwdZrcUP8twBUyF6epPyJrc4b2vTjQ+mwWd1xoCQg8BF9ts02YTecx8A
4Sqyx0d0mEwtpmJZqSku0WvaEqoWaOxabU9CINVu9ZUJsudAiW7zFgbXAdVfQriGsOVWYKKRwoRA
fcVdHE3R+HBrl6PbfsW0V3+eBfRLpvLjRBXEBDp9FVF2KjPHojac4MuFlif6LGfs2F7S1GcwbR+Y
y42uW3xthosjHW2htg8CqJiG1lKEOd4VVjREpztu1Rs7CPRNHg8FAowmNlDb0uGR4FBs/eNUhx4D
9pXtYrK6b4KTFA9WM7ltGwIjR2Vqj+oY+c5i53CHgQ+mPu6efWaDDCzvM/dXwdEbjul/Dg4BWXi4
BxjEz3nkKETuzEh66AkFc2maVbe3ch0Wnshcdt4WF8nfwE+I6WrAq866y8w0RArgKryIHloVf9FD
YHOFTSkePJnoEOtJrZyHo+7z6XWEUQFZ2ikMAJNyvp7qLvlzZ86BgJnM09+TyKu6Xa65Jq34a/Lo
mE/Aj1YtaeVwpL8yDUmp5tn3FaCLLebes7kmulB3TV1Wk70UDrZydCXg5f91SiE5VZU3gQ2/oQRA
YGrIuZhzLsF3WIts2O4NMIzUCJLcHI/ynzeWq2C5uA5f3aAj/2rRorGXUi+zxTxXVlsAyN4dRjfw
hfSQ6t0ah7ihNlHEg3qJ8sscP2ttvT2kTRqJpXVKKoIaWF4iGLG0xHAws4RVXu/dW5eKWiZEWdKH
axLNfVsJtLqhZn36V+DQbR9A7jsU723qZEYC9ZW/7GBdNViBMiVC2H67id2ZfNtsT0AR/Rwuok8C
HP3QqQrgwFq4Ch/8ijEHymTi4kSSujYqauWjxRaNxn3FPYpq8i7RkhGVnHIIhAZzLan81TwGKIfR
2UU1ATJOS4tii1E8Z849eYv6WM9oDObVi8jKAdHLuuhbiTZm/0PzumeI9Py0ReSz0d15bzX2R/MT
bE3LZfPrMWQlW/oTlXUS+ur4tKL4zEisMHcrOgue5FabUV7t9FI50WpBhm70zFaUclXb/8yE/tJm
by885aFiMcGf+hFR2pcW5cXma14HYCOYGrfCc5fGoBh+XG5rOIYb8uCvIl/b8CqQiKcL9DU/b+br
mYJOyl58Z7CzOlVkxSe3bRIF+J4MmaRZe5aNejSznuPl3fAxTG4ti7DD+Id/qXWWxmpABQ2Wdyra
P4Dgvq7sg/LY4Sb4qUEi2GTFBoF4/Hz7J1gV+O3n5D/apzac0Epkab7ZIWbhIWoctaYzuNDQqrlC
EI/jWGnb7gSOUo8NlJs0bmMQuKdy+kiNNB36h5VfOiuKP3ApmBi4wd/S0g9Vk96kPryqrgUkDoGW
El7wHHU/56JM5PxDzlLlh8M/wJqRRbMudnUSUxO1jGxfguRcpop8OTfJQ9JPHaT3oice7aWcasCJ
FaMlI6tVpZIFTjm5hp5dBDBeC9E/7/txA6Ikh2+Hx8O3GagKSDkaFYeP6NpcmJtcQxyMDaIaM1od
3H5Ph9FiwWp284m24O1BRD71sGVvHodi31ANqj25y/fSLp/H2x/KHJtIRbLBPgvnCQf1aiqCeIk7
IFBJmcnT9FSfVF25AZOgHJIWO/4kSuSPnC4JGopl+zqjT5a2Mdbe3L+QPMvc5rZ9OAbD5Hp2cPGO
zja95+K0d46lghMGY+/OYa99Bm3VCZUUQ64H7CZHL+WLW9KL8LiHVBn5R+tlvIjQJnkH1tzuCSNT
tWMNxywSIKf0+fTjc438qtmBz3wY/MiOl0w21nYgM8Jb2QFdAcCejSffjsUTSpGD5W9bA1hbYrGz
9y8EqYfaxBdZjnI47IXZcYvbRRwDm9tvT538OnaqiLJm8OcZx4d24OLDvw41mVCPUP3BshTKOs1E
zw1l9hlByuz3n+RpYuKKknpdpG0qzpff3IwE2k46jyR9ih1Wh8ZShmfp11ajlS1uXhJY2RMNv6Dx
86/urdsDg12NyXfG+/LGvVKDaFji5XLGVxF4zbybTU7At8x+6gmbCOpuwgD3+2FpFpnmp888S9kC
tg29jjDaL7SdUhgV+5D3ePpH07TvybVkhgKfNkAcmRM8MpJHpeoxn2vksOVdNt68LT/l6nuaMksl
+CyhCHcUplBqMJD3jVIpSASUgrR5ResXC+jUjZFn33quNZC8cErAPpl9e/qvLzgNpXCI2iXiCW09
B82zpvUAhoOgFf5q5x+oFovPoL1P6IHdAhhWKmTOo3GUztzs93yQRglES8C11MKyaDSYlsadaNfl
YRXPIj3yo8bV23dEF/Vm/Caq8dZwCodQPtPxZvx2ZaW9vSQ3NhnBqAUQEq9yOoX/R6qQhXhsBlJl
RhRBIXPRJc2FgiLHprs4+P5UC3HAYOg/GnULFUEoKf/k4rptF5xkXkt+OR8Fk5pGnDZYwvUJZfUx
RSIN2xRdhJuplgdIURSUME6DXoFj742H5n12zyHu2ukxU4DiJsdIurBRK89sFQtC66d7OOd874yb
8+Yd1KiOO7imn402GkUiqT+7N9cYlbzc00tCQoJUKFis0CQUaCaxp11pU0ztl45GFPoMXlaeILjL
Wqyg7tAajczE9YfZm47uPtbAdgvSnFibwt3F0iVFdTdZplmfxHx8g8wO+wlBvOm/AiTkl38Dcsg0
+coLTeu39SG1fmGepVFu0Z8GUhhB9EsOVZwNfM2uoRU7OwwW94VZy8VtO1g0NgYsznSaifS/mPVe
Jnf/+hoEPqUWWfbF0UayMGrkiDH9cKeRtPpw7pG/sy1oP8t0u0i1irY1QmLheGGzehXhFK4USBUP
vCYjsasYHhp8sxXvG3ObzizTNDXyIO4c0391/XGN949CHaQqBTFgAGWZs3FQFrA7BpAotX4rUnLH
qSBewyHECIiSd90gmhgcyAUl+x5c1GdJRvUynV05aKWo0WmGiEqQFpMFmZpho94QCrK0OutVPh65
Pm/r35raPmnxnsMWE7os/b95FndmcSU8z6X/xxZ4dyXCgJEPD7lUGIuGah4kNKM1u0gereg1UZQs
iQSbNxt/lROT9jC9fu/Nn6FlDv/WZfk0Tuo1k7SeFBmF9Rn8MGLCMo5D2SVvf4DemeZjeuR7TaBY
hwPz2aTBzu3wfWBsEAplGuYUddTNpwGEpvSBfiaexNw3ifjlNedFvdKeW+ktXED6i95ZZl72UnhW
UudNp2nVVIc58h38CKGtrSawDZTYd5ijF7Wn/IKEAw1cnHA+ukf4pW0qQRRCJwgxF0el2uiQNz5o
Lm6hAzZyPISR2gbbe6hu45d7511l619RoSqrmp5RROKAKo5ZndA/yyr0FD42ZHACLmA5jHnwxdcV
Krx50Mp9BoxjijuqO/TOqF7CsU+Tks56BLM3OTzoSfdNu++M4mAwfSLZinjyDKRagLulyDotZzsl
1hvGqrZdi+XF8SOA2aW1mztGgaDUOusqgRFYc8CZODcg8UFygDwy5emQhBbkxSHRWF1DAFrRQQPW
mgriiQ9q99n2fdE+LnHqVZxnRoilQYC2mwpRQVUT5nQ13PtEtPyQqPkUOkOzCXtMyfvi3nEus3fI
r3eJveqZXpLwoEzko6ez0DmYpaxnYHunijnKyf9HaKI0Klzn2YGUc1Rxe2bFXDIF+KcdFjVRx4UC
+uXqovZLr9Dzg7zTzBFnSr0zGwftMaNG6DY6e8k33xtLybJyx61OX1IYvkBEjIe3qUDkhiUu14hs
tgMvpjK0p9vXm0ZdDF94nwdbymOFD04i4sSq5UbBdNZ+BAxXFc103NrablWcnDNjF/PoLuHxQg==
`protect end_protected
