-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Y27WD6jjWSQzd3NkolSUycCK2AQQOHgI23m9SduGqiYJC1fV+jer+6/EbghciWd17A6HON10LI/D
9mZSZzbJxn5MfONfOuUX8tHquapypTcGSAInsp0vxcp1pulQHarqSNzoOYQbS7gouFzcqN75/cIn
/BwWGsCVVEBfLS/BbU3WLdT+CLR2sgYMR+jqWjjZaprnpoqQjTlaCo+W+0k7tJlcHeWLUSn+o09e
6tjI8mRvs4nWOJlfyMTrlGPE3cg1FBr7LjZigXunrpbtUyxpw2/pMdfpUvpmuaPyvRNRQj4oSMYV
FzuUrbaSC5CrVNDYggQWPr4cOLF8D28PEb53IQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17600)
`protect data_block
/AZ5++1f2+JbYD5JTF0MEurg1OpWQNEn6gy8BZ/mPfGkwbGEBrittVd2ushhKXqr2zE4xmPgDCbJ
T//lUOBZijL/icdvkhlpX8PqCsMA3eDpCglvmSksVXk2yFjf6Dl00OAtPmWuAsFcZeKbOsBwS5LR
RZB2+/lK0mjWmb+8CCbzli9wdPsqg22g25pFCPPGjjmcbBbJY9i3sQqDt5uTTjjDzUC3vjMvfwWW
NkhV7Iu2EXDJnRTR1VYUd1asRBlTfir8SiWztDN03jwTgXZwZUyO/ch47c9IWwh2NQh5ME8qNoJx
ZH0nD9vvXGXeF6LQTm9h9bl4ijBqyHh4QYiYqq54NgT1R3wbvlYHwvm9hsnZrV0RQqpbdCkNszdL
fI5GwH5Z4YHXxxb6vAU1JFf23qdYo5Sx7DwSKWu/4cl9OXnw4+mdMSRB5iQJAiPSrMAjBVOLuoEs
nMPhcFP+6FbjJxxX6R2xs6ArLPWHdqX5UbLdS7nX+gdA8oCxQ6WtipjXB33pssvzj2/dL2zZ+SW/
yxKvxBC8CG/KmjSI1mGmuqQ+cYnhOSWeDVe5xa3yMEsMkNIOHrn/SEFAYvMFGiBO6fxtSuSP1xmZ
ldHU2xhAofuZOTQbp5Eswl0WFMLovaUfDrIi9/GArGMVPqLcjr9jvZB/GLcMCERcxBJutuuwyj6w
tI8hQHjZnLq4OX+zI9WS9eEyWTF9fYfan+QX2x0yTv7mKMbQ5V9VMrAoe4xyztW8t3PxOOTLQOqn
/eLlHEJREoJKnTJIX2nBJ5DgmIkX3WPDOVwTb0jNaQ60pLwTBMKh6BNoRb7un3N+IqvDxaHMgnRg
yJxs1q8gWgyTG4nCf/+a4a7kOJhRMMsohxZGm2k0c/KAYIoBH6YEcOSDiH8yM2v/PBJHU4p6Bphs
ToiIxEa9T7lyJrkbyuSc/n2mfzJ+UMRwCxvaqAQJLk37njjR3KZ1D/+nMJXwZppV5W5AZ47jBoA1
xJsMYDtvzclTpdQ0Elq3oz4mGyHOq8G7tZRRmCrLrHGO+khSiQ7h6t6q9SSikFzhyPPO0qwE5i7U
FFx2rGttiAQG/6eWvxV+QULRp3DXFY31RA3WdCL+yAs7brz3cfaQXaR3jdKuX09QjxW0iIOkTXaA
waL/BMkINvY7N+f11rP0h3h982IKaUYGl6VbltrgJh0crmF97MCvdDIEosOvp9Y4Vywi59Nsmu5S
pHlL/JaXhkDYkSD0/T1/i8FHmtmNPOafkvOZN1gySFZOUrz9bBgoPQR8OOH4cuO1fWyNEX1S0Jcn
mVaVkoJA4if2wO/1CFVRDtQ/rqllaMd+vQAXFCycP7AtVAeyn1Z354JyCkI5Xr+GLYJlkB2t14la
4btoiXpiFmX9TVgfZOgWk6pRXXUYghdkdQ+9OTPgUlLDG9PlzciIGfdBMywIK6Njnm8gmLiRFoyA
AdpkdmBNG1cFEstqxisAWCVALVhcpZflS5U6Lbe0g2RGNc6doU9XGBT+lZE4GvjiO70nUqz1NxR/
YVLL0dAOek9e1PlMmE/tJQtY7zn/cTW0fzw4eVPkOdKWJfb+qb9kA6pdchtB5fzZ4Ggn3l37i3Cf
0IBGvdM/0KwDjE88FBTTQgt2FP8dl+dmSu4bFxaviO10z9VdPEVRxAszraUOekB2Eca0PW6qZYor
uMVbY1qqZJk6UkjR9iP+XSMhmlOlRgSYuwkpfZ1fvzslk/Tx+pO/dUKHNmr0Ua+vM+9cxjSPYkY0
FubZc6TTxn7MaF/n8DTxCF9F9EOaxupl031CVFGhsQOW5+ep9Q8/uCbvzSYkVuzdrzk9tHvex+Jz
hLFpHg96rW4aVSVZBD9ZbxInhhEO8nchOJoqw69GxEyS/Ne1GbjtRHKBEzoOGwwUENsLTDMERrGr
098uFjVRPQzRLVLeZjyCV2fwILZIINiSMfBeiU1cBd9Vv3H7kn9YcvO+xvhS12qdmpPyHmtAEvHL
okvWo9Whg7ngwVbzgtUL5oinaSwIOW7AEVtquHRjkzRfsPUEGi8Xf5gljDcV9xtjrtKW5K/Q1GLm
8ctkh+ENgXyQEIgQ0PruBQJLH5j/89EeMzkLFvbUDRNUT+lzVypoHu0YtZkij4SObhW1A3K+DZit
wfagHYrM2xMYuAHxIN0sp6A2cVxSbPzBMm1ALVDJ0n+/S/IYDA0gmj58o0I3yqk2LeLhWy0HiAB+
6amkbWc//cIp6iOztgs+rAnuNhi7uE66D0Pl2LJz7ezK5txISt5Nr/VvP2MAMt+tsEFcp4oqvkml
taT2hAzZXHEK1OzAJYis4aNCtDfbTEjDhpZaLfILsf5j5a1hhMGwoCbCkEuVVXlUjy9n7ds8zoAR
UcdbPRW6ogro8PM/STjNII8YOBL38G2dqOr54SGZqu0LF6JSP6xLar3gZexmUYw6k+yApfRD91xK
Aog8ktWrIx3X98hPYQ+3cEVhP9XgLKXOZMHhuWwdLvAkDd4/sfBsbTFSxQF3i05QVA1Qan0hijED
IoZ+GZSOUo+maII+EBPciuN6OdHozq6Q+xeXSXDVrfpZFOUN59w0BThyE0WNWS/6Lt/T3gfio56G
6x380G35y2qX1D9o4LFHCnKYguhWNA/edDqgF7jRkKXESKkb6CNR6z2j9ZFsRIsOtLwUiGlHn2UP
cBmR2OJq3qhwJMYqGOwP4uUWVJU8prK//YlhFgMvIrE4FIrK8QXyXqf7UHn6nmmSld8Ma7oaICqQ
PTjCVuWL+7YGy6z9tpKqNAVauoky1hvE9R1xmnAedbo9s08uESfSOQoxqY/nuftqDHuu+ORmdrGN
qHmWnXd02Z0WraRzra0lcFx1+EXzqVexpi2HA1mByxQwSHeo3GiYyB3ZZ5YB7O5SpDTB9ErIknPO
E2c5muvFtskfg2A7uh4960cXO477jdpEHG2kP9uhCVecNUD8VfzwF+VSAQAfCd22V4xK8wPXEYNu
8kqF8mWO3V8mG/jg6FBwiK7btfCiWtTECKSZEVqIsEws+9cY/zlv1HFQCb9HoLusOWhqmQwkV0vF
SvBEfkYF0pfDrducVBHDps03OEiYpziE/eP+vD8SC1bIJqR4CE+tZ8seyY31hvHjPEGQcPfIO4Fk
mFJAbg7ak+miMDlYNcUSQ2vP+FH97wh/5J+Jokd8KCiTmJ/KbSNK5zBHYmVoNo0KrmSE9W4k4ABq
BPdbYJyuxhes0jqiMWgPsNgpwat7LMd62w1EpyUw9KfvFtQxMSFXqlwKTFaD5U4HRNYp/rKe/kGM
C3+qS7rv1a+Ue6ylzY5QFji0dEx/6CiXsOTOXCvZgQRAJNLnCwl+/pwYPsCxD0WfBuBoc54podYw
XBh1cAARNv6miT2ttPSGyZFjnJO6rrK4DOz1mE7PExxWS3FmxCLFM6QKDlyGJTJ7Ru4qoP8Un8ET
J6Asf879Dam8k/VmUb84sWiLhzQOWv0xdKDKsOw+W2X6LNE8O7tZH4mhXgu1D1YsMXUfHwqsbkzD
ngzwXSQH9M2MfGmVpEPVxN4pdbZp4SuJCfYm34xjlD9lFUGhufH6uujm/6mJoov1dywl3i35O20n
ABDA15BrlASY2c740vqa+qhodJo3EOOUwo+8AaYQ+cZHG0Hd/fFvQK4+kjMO7ioeIYZZkhGGKHmz
a1C3EMWbvyW+vowcuV1p0DZS3urJ3KRYkw7ocsblopkImGsLKYjnT3nq2m60gOuZX145+eGk3Wcc
Dl9ZXaZgiGZ2BcgGyphYN7SR5TXvNIXZgnoQ1kXlSEfdNztjYDXrymMCvOxxGlVfRra1JW9hNQf0
JukOzXEgHtqSBzq7WbHtnsmkOL/ZjgFl+ETCdHb2uRoS99WaSHmWJEJZEtRwsY3+KdpdQ8QXNp/1
LgIFMGnn0VMme8+gIeHo5lq34XMCG8zSe6L4RhsjfLKEYjMzEVp1dXz3D/1XG6a3PArsTWdobgeQ
eqs/Ed218PagmACOD//WwhijLQ1fsI2FYYHp0Qu7EEt56xG3YUTNfALVHF8+BbSU77DDnZpziDbk
e7SyA7gl6i1OJqdL09qFB82WzsyG4zy59lrKlvkdQXLwY/0t/h9v65LrutNJGl0CrErmydw6etKu
AMVSbta2a/jfmhy+eDmAHoXQ1I0UPHBn7vlyexF742Stt0oSHDLXvtFLCNXVBVZ+/M+VSlsTQhTv
3mGMkjPNaj2AoG75/Q/YZYzFDuTq2394v1/v9gtsbMOK6oUkPo72w8z6FnCk+5xB397iQuTPdLdv
U+9kXIy8QZGz8JjkQYYgAP0dhndktWmD8wiVrtpZnFVtLmTMgfHWU8MSpvQYEpyMFMv1edhCxIEL
LCcjRJSlToRgOU7zcMqAgn7S/FK3PJHc3VmY5C61mTKoShEOUsnr/QG8Skkiin/S6vQoeql4DNSo
zLGuFdac/XzcckJm0cnAgsvSyYwsrnhuqMIEdiojHjon4U5hQCiBRTgSsoBr3sNVfi8JdRku4I1w
f+CFYaFtHv7RUebNgXH6zvBD1uJM5tYtH8VwpvcJ9ukrneCk1Ss/T+rM2LZDEAdgw/J+f3wYYXlQ
cZhEq7Du6fBS6wxstAwDCbSCkatdl+awsoBLDwtSw6EVKLeJZ2rHOtU/4tes1nDQ/mQvouUoXVto
/1avc7USmn5saHpGQOaDrcwHja8aMdtSDkSBevO1gla+4dhXkotCOHRZy9oAFMISLJWcarw6jbXs
TCKYTl76E7b3zz5UnMOSWhfWYwHJ+Xga/r5KhW975PNgHbHwoZc5+Y0n1ZJKbRen8Zx1DU0EDysT
UaXue8u0CRZ9nVRWD33jpPLi8CTDFCv/mDCJszeaUzQsR1WmkgwbL1YllTvnFHgOshrL9j96N5Je
rp+i16RSs+yPXh7KJmFbnk9wcimxzQFafFQCfTTvioMprDcj+keQl43yNBGdsq3L/MG5OA+5WI/7
6DK+m40NLtJJDtksjn6aWIIMER/4xoKMOj67oJWtqbW+fh3xeRaWo08NC6U+vvydyczZDfjkXn5k
Gt234yU8fmkYwZ15UBrfKmQC0vinf8QEmMM4uzqt83J7ufXrA+a0R4R72+gOXsHCXXLG5mUfqnRk
grNZ3cmFnD+HjMlQodqzwjQfZdKHkqwjoMXJMiv+0spPrA6MoZtQT3BM15Ocq2CFuVUC3jK8w+mH
Jx0xclG8e3SRMlsldt6dbMB6riHFYDzK7lIPGWomH8JDZHWMFvepjxjVWigaUs7ynPbdsluO7C/4
+TQ9Uf/lU9Z9dMT2SX+ancPGQ2xSYEynLIDg+fOXCqWSbwuk5xnHu9am+ewcyGN/aPh9oPRBiiFc
FOtfxAj0kN39rXQbY0Aztj4mmDt08cDamKpagWCO95T0x2qHVOcO2DPsV/B2ZX2Vh2ZbmNDL9Ilt
wpdnVkLGQmzgV4O8ZpmqznDXMqNyjS1O7eCTA7cMEN3cKeH8Uqp8QLKpQkS6DQ1BM8ih4uzkpgga
lnm4l6rWWiFMMqAIQ6LE2MRA6DU2jJb9EaB8sC6m3/fXywrGmY96C4f1woDx6NB6HLDQONDa2TfO
lwJtpPO1Q4QbRRJ6DLeTKZdnrgJvN2/FKTr+lpgBNbaB/fT6edGXOD+bdLQY8UpJrI1n6y5SrPZg
7bM4sCvxF02ObawhruDXEgnrDaVU+d7dANFKX6JXsM+JMlwA5H3cHKMaKcGqtW/VW9YrSiWKw/Rj
9Dy3AaKAxvzWZCt1eBdvpfoH3Kp9askzLrjQkpa3mZNN+vIxURp7CMtujra22aYU2ZidmiIZe8gx
HXyClWLFi9q2tLmvOZJAl1bmIaJ/cnYmSl/AppXs5wDDHt/q0mGm/eulx6t9o36I9W4zRr3DNOhi
JLjswHmsMhFPXRASlVp5DU75oZpfAQ27Vo0MnxxdXGBBOIQgmF7lVr+iCYXoL8BSwaB3zDP7IQ8Y
dEUdkPzN6HIRxqdWfGCQZebHvoFKomZfbivJMjB7AnM8rSFC60rhVZr60WBqh1o7b9WKarSrBRGn
+d7jYSX2sUod/jyhyysoU0UmFeIeFuuZ2jfvPCO0BmrrFS8x2z4AaiCN5vYSSmykGLElgWNELVQa
mhM1QLhenvkcY1ZvEtrTcErjBwnCGKLcHGQOGCapLzqkMQWa52WQEuHQrCBITF5dbzeH+z2zyp0O
wluF/SDVG6ihUCeKapSLw43amcO+a589WI6D4G3IIpSiG8hQwjmOgkp6Ie0NOGw1d4tO8VGKVEzm
aSvNFiTrIUO0fcwvvP6q3wiAnw3wCmVv5+9kl9Qf9xI7GpOi8Qf6v9WIdavUhVt2wTkg+jXdfIku
e5uWlS/vkglD8tQLFdBVyCI9ol3yUqBym8rBAJbJnx4JQQ22nQMGp3AJjLF2f2uO5Nikecpn4kV8
qpDKEnV5zDqOfk4fTQq/jw2jnQdx2JtGwGzeZQrOATQ1dUpu0DM7zvcLpxXiRpk5DZ/X5yULeVGc
pLaomrGGKJTEU/TYsTjE1+AzIsUvobOs49tDgo9aQzzUqaYQqbc3psyTRTqlianjizlsPqMsZhDd
lE4clAlsKUi5kSztePJdpx8KZYADMP8qDqSwT1h+BdUpA4jFLN5QSSELbHE8E6/73WIgGO2GOUAf
psdsRF4gBepC11fekb1xvTQeewmou50fbrQSzBTblyr76apCwZe8MKAQiXbyY6PNZmg/lcy5dN0B
yN8I6LmclPO2wZgRRzTjAyJsc+Rcg/8wCj7zHFdk5JLNLX8vx99FKfhVK41ZYroBbRVzX0UFXNws
eBDvyX1NrZFS3JjcyeJxcIlWT9pc6owaEUYADtmb6yn2aHBcdMB6HhuNUna9Vc1cnOYHwcUI6J8T
BjzirIDmym+YL1Pho7iXXuX5hZRT/Z4/u9gHohS2S8n4XExbt6HyrFTAgwBgzUUwgPXAK8DDio7x
qnCsi7mtrbR/JVztkL5n5SEBsUP/2y/C6gifGUcCzoqtTfGR3eT/XmLmXR88sK56dhZcBhPpdR0j
CWeK3NPEx22FR1Lx8nCYqGp+eogiQUmN9LlQU16B63oiVBHAbr95q7KIuu4L+CPQpdvt0At3N0E4
UaQpjVx6N0xUYdlYz693+7Qn2N936fU4YUknfWs5JtxncLPAP1rV1D/uNLRf/0Pu4uc3Vd+vVDCZ
h1I6JEEZQR6bX3Okec/et5jAAFxQmKlqTsMtKd0fziHMKSJCiAs1GT4AWLYjkDyVX2KcQ1YCXNbM
O69ft7WMJyOfLsEBN9y8pSxrMvmJAr/aKhwMhhLa85LuQkPJyDb53IEkm+Vbh2EzuBNTuG0zJk15
G8y83unZiZJo1nK5/6l/WrAVFf3D5KcvQeZ4nTPn/VaLMHW/j3mPZyECPCSWgQjH/WoUSKMfHQjJ
qdpFeXi6mc8ZM8qyVeqMiTWJFJRq1GerDNWmySmEI+7lprIA3fKqmojOMAnAB0RnYEp9SR6F99Pu
0EQQ5rMOQDKmj8QUG4fg5sDt0xtyu1QY8aFer3ovarZRoCGTUQpHrC9VEmoJgk9mAg12/Rz8kUKi
IrPAe+i9XFms1O7b/yZOY08pKdcPT3UhmBH+pxIqvNaZafH2plqhhL7cw90MzR0LVM3G86ZKVKTN
vG8Z9araCeULyCudFLaKoJSm9SeobudN3vvxspkd7VhGcRRtnWuckHghu5vR0wXjT4ts5r3dOnGh
6UZz3ZnN6enoo+3mGmhK+6EkGKSSrBuW9f8dxovzhOFIbLYyJaMO+pBnax3gJVK32D/Q8wVesDu3
w76cfCXz7KbVGGBbnjp3ppX5sTxxqYLrhsX4P7P8Afra2bCpdobazx0zkhIq1Qt8Cu8xZHdjNBs9
HZ4YzEPK9j8osL+d944Koc3/WqHh/nzAY/oQRazFcoLp8/NKJB3ZyWuB0e8KciUtoGGJItB7b6Yo
s2PF3f7XfoclygfPxHsvYlREU12u76Ua/p5YXP55HyplOQMiDBXzN1bVrK5/fxC7efyLeRU6i1rU
m7eymNQ9DgyjuzNvzHebAUITiEN0PD87xQG/RJuHPEzMHTmg7S0d6Ia7e6nB7UJ65wRxQ/vIGeP3
VnDm49ignf7lfg7adQcwYy+xmheNozPaocHFfJ2jFAYEHjsfZQ8FlcygfKe0EUypF7A11c072wUG
wWDGr6SQ6gsEFRiCNpJaq9enViGOwi0WjvYqyJRP+so1RYir5Siyt433wlMbisWKur6ync0A4Mzi
ly7UKD+QEXABMq6F3/OIEH017IGF4cyKmyhFPsxP5d9xj8wShss/D/BFyqFiu66VvuNK8syoZ8SJ
GYDUIKDo8PGaAv4h8FE4t9DE+J67pagapPsaHrNZm+0rSiiRY3rO8id5/GjkJHMqymBAAHbxvivy
7zY6t7igltJC4KEkw43ScRmLaK/39lvzh0x5pjvIt2tcC3NLrxNpK/Rs507Hbr6+zayobidVboeC
Ju1vmt1dZpUcDB4pQZNeGYm8ct3a7Hy9BbBZes1bRA3QV+b8FmouBv7Eb3UD41DPPO70STLy5loW
VJr5SLedqHBxx/TnQ1qhfn/zBmfn+kgVPukL1gSykDaAb0HAFGxpgxqeGKLN1oOgXYl3D7rN/ENU
rTRTdtxlbrd4mQ3JB3E8O+dPHfxYyuwLWFtcQWQQPun2pfPb5yYGW/StjBVNLjigVT8KTL3BA4Q/
cxbXkuCL/IgEA8cwQu6gnVwiCg/n9701dvu7sj49kevfXR06UBMStbN8f3u3vJl+bktKa1UWO/fY
wvZs0s5HKcinqA5v4vXV7bvb69mVVQBcTa67vS94Vz3C1/yGqMOiwgQ9XuzC2jnT7hIovrq8tbM2
3LyD77ehHwN3rix2J8H9suj3a6K1cyc5awuUjILURlM6eI7MFtEt1zFvVoyuT44D0ZZlplFGqqBk
nptNStY++yDTZLhoGtWu6KJw3darKlr+XvZX1TkMYMjZQcH94+Z0gLFPYy1hx3td6cINACut8Ghy
IGns8y50jQeLOcORU+2e6oenh/JZ3hKPGVeNBgxG/yr2eornlharO/iWDAVkp8MjuIvP0eXNOqhz
Jmc8BXnYyqs9yaZ+wcE7NJXifXhl2SVVub0nW15KbgijYQUbN0XQMtbQ1YYFHYZBYwBnaVKFrnjd
i7+FfbA3C/UACU9ld6ZlbRI3MkQBGGTOTNZ0lW4CoGCRljS69ipbQA8PrYrRZriddNhDedC+Qxb0
w9+xSX+cWnGfjtakhco+Tiun8MR2T1GP8fIVUvCMmTJrQ5yNkGf8a4iftWlHhCZY6wZMdBEdfwAJ
EeMCq7aTjQN8gmMpLJXaaN/fNqD5+VG0GaDW6dvEjBn3xdJnpCkSU7vWKGAiG6ptHoHpp8/EuSLi
h/EA634VmefM/RGTzYFXYOSRECSX/ZL3Nnka93lz8mWzMkQyqQvffAFgEgvItRO0IQT7LFenAahv
2XIBPjDvPgpmoOsxRNI1V7eXiBmocJt0iwY7aApUdh0aBD8JiuG3vOvPpQlckbc9e77N1zZqHgJw
A8T0d+LXG2XhFmySYJ5h+7qLSQDqv2M11KmFAeSu33vm/6YTsM1ddaHY6V++c/ukgQWrHFYpNbTs
IJyD9+wrAar1VjvTqhL5CnNGfH3PYLYHwDOyiujnjARDEOeT+CLm9fBfchCLYR1/YYOREFZhpnRa
WKPjKPWlbcoWWBGBRKaKgVovYLtwg4W9SAipUeC9dUDaYbEiS704oFfPB1wr8MpTfFcelzoO+cRt
FJnC167xYbx+M2EY3lafMhHDJOnPR6WOl061H8HtWwaEYuWEvxaJAk27LnO1S8Yl2Jq+cB+K05VZ
ob+GU53ApiPAM9RmNk2Rfr/xeQt5Klir0SmpAVAabymJv/6ViPLQAfGXb1kIJU3AwK77YEHRB4MT
WoZb1ZsZXIZJcybhT5QwoXEfr/JJTpqF5gDjEo4Th4XSihXzp0AYIX7RGz1dGCOP/mcgCDNji6Ai
dh0hkPZzAOlB9wrhm0sTIP1dne1tjVL5vGpWJWlJCc21/ho0wd+4GPNvsXEh5ANaIywZ1ATXe5Fk
ryRczxQB2gGUYpmlR1DYdKgO7HH5WGXNV9aSahXepmYr/Qo85Z7SHC2YnmNrgt4UhRrzvM5vDVQy
9fH7qsjJ/jazBSdgaX/07YAdI36/CsigEf0ltzozQNqDfb7lt8l93udqBDn4vTLdEE/fSkNYJIxp
N+npe5JyDGeC1oMiqP2P89WKEdFa/f5aCrpublEKjHcF5YdHlQuTAeR8AkACFSOmIEHSAKdNnlvZ
ekJjhVQMKC8g8dvDrwS7U+LJC7CeUJqE+64S9pVZB0ADmhVPwZBdyO2HrSX99cT2WT/ov3QeGPc+
9z9wZ3o1tSIdvkOA7IPPA5U7FHzpqrvOPxaorbfN2TBN5OEsVfBhzrJiP+/EzVTm0BKTkdR6Ul37
SjvLaFz3Uo0f3uhqxcpgB9SSjYKRMHQi+ijLxGfW7oHpL+/9s0DFytZ8FcuGqV8PBpdu5MVm3K/R
9Q6I9jNVz7uysGPi8jMAhJc58RdgA8xCDI/F24RAtvUPkKxtlXi3iggElrCbvUENpNs531KT/ZnV
dahLi/tTtHGP4MSbZv3W/9woewDf1Z4gnpqWcoS+hnnakHH3ukXUJ7qkSFlR5aYLBqdlEP4XTrzA
AxFKUa6pybL2+RqDz+z0Q600DI8jX7c2pBJvundzPe5rCqVkJ7hTzeNW9MqgKN4C20bq/qemCm1m
UlMKkGl1PH1umHOtkMIT0UAOH7vBEwwJwSedgnCw7fwzWkKaQAIZh/DEgUcMder+qbX0WeXey5YC
5yGLYO5kGqzPGvbwd5y6ZbQiJKdZctq0OmdRECZkh2zNLH8CMpTSS+DTG8e4DTBq+jUjNUnoI8VQ
Qmmvot8JVvHl4Rna1brHcBxeVv6W8Om67IQLjz3GIagDHchCRGzTBF49QgQ8WbxlfqzpjFNE5SkA
3VPQYKiGccDTOrvFnbcTALaZ1ZzgkCW68Egp4/G/vDtLKbnbStyvaXJ80U8xnt9GgIvqrp+TaW5V
xHHcpZjNmL3TI1SbL78fcuv7p0iamufmAD333KdiDKLZFFZTRV6r9u3iympf4Ruvzgm//9ZNY+l6
mN1f4tJBTHZOjeI67zi9gbYP9nGj9PR4cYQFekT4VnLajeCgKw14NnZytulzwmYc70Tfnhkcibb6
oAZID6NaLkGhtTNukf/feKP8oyL9f89d0VL7r+ufpRweAxwexoWjCd5+YuM9u4QJ/qJzfzWk3UzS
S7wqEZjcj2OI1279ESAE4AUOCH8Gwy0qX4qSYC+Exox6tdmd9jDQ6PgcSRW3CHVObcti5PnJcrKf
GeaiW8AB4an1ZDuCzVSuMmxyxVJ6mIwqbnzYAiVlZUdOUfMg2SgZISe/Tz7S/vaic90+RtFhLaKg
x4cVr5ujWYk3OJtNqdV6Zn+4+H/WQcZS3WvqAgKPf5/wzOdhgyowPYIWyVVelcmwgP/mni03HarG
KPqZAMtLqhyOJUPjTVY6BqSmBNvDjP2Bal2JtKgQAfsHepDdxBdNE2JVbUjNg3EkJRHwvr20mE2x
UdwgvClkDrNZ2oD+F/hoEVWko1+ZnzMOeoRTyysJd53XgEXLEEr5Grahjmb01KTNGzEjffzyKFv1
CGQK3Dzq+475/QvYOGS660dHJ+ILx8nYkH6D9tzN6szYPMsUkIIrKPupt/2BCgBQqwISoZ9TG89d
IPI/5lez+oZi3KSfVpfIqVHPzDMymXlJULuefo+ly5eI3bSYDHAs8343C9xFNRJNZ7dnfPyW1yWG
Z9k8PzCs6Tbe+8fQOzifVjQNr2Otezdfg/VgNW8Fa+SFmrbQWKgkRRwy5HCno/GPmUT58t8ZEpe9
GokPIk9vomfTx9GDMIWVTXmAlI7wW+6JfK/gvCrwnT0c/1XeiNvEvK578Y6UbtyzCeIBDDoFso26
cmnIFMn9Dzw1hhGUwmv8eKUfT0+Nww4Iu3Ihmxoq3ESj4XYxC2lfLh6Yhvm7ox1psPGTbnVG4Ci6
uU1gSYz1KZ0aAEnfPPbN3tRvBSrsvAoY2C+KdYtjsZ6ictfnV+nmUfOLS2lR2xv2P7bJMHR+ekGS
pJ9icYOuCTFgYjxDqBFhELz/O2qKlnX2L0H+kBlHWNLRD0ZCQ56HISCGuuoAwWHjznPuEiefzAxG
7Zw4ZEbYso/HGdL1Ic3FtsQh0kaJkEYOGSUMJbv4S/iezfpoLJAyTPcRXipyqQzRQMsXN47CHKRR
RrLAEnbf5FZ0XvSjGpSskyuFdvXRRCSMoep75l1qk5eoCLhnZbYrZGngJBTcdj2y3d4erajxNd73
H+63wo2ei6/PGM56MmXPEHZ9BQLRj314tKEc69umaGKVWPIH+iQnY1GD+ifMqzYYsK6YwbfJ/FWZ
m7ecvSGTjndXc4vHCYsJJsns00B1rtajaJgrERsm77KAmKjZ7KKR2pzWTmBYar/rNiLnsUK+wjMv
80+7A1toDPzNLKrhhDNn15BX26wHBqArhplqU2Il7QreC5Nif0pZE+8nuIlCl2GODAP6kNIBxuns
4FH1T698sTAPmV+wJyOv5Pm7UY7mMwl4M4rX/T/au718xdVrlLtuB360/9pi/VIYQ/e5IU0EFYUf
NqXGs6Movlr3I0O0G5lXKhUVx4rixmWhoRC4tTaJMjNpYa9LuIo6uM/ObykA8QDbfl86PBieU1B9
m6hFJ24WuHsnDamrSNHe/e4sD3C/8ZyuFwsuSRLIqIhDQ8luMqDIv2JbH25KTUEel8zj6y0WCb6g
0/eMOQ3Pz3sEZ63i1PpO6Il5zkZuLmUhcWkcAKwV6uSHbt6nwriqurX4SsWmONQ9tpj+ydFuZA+w
N0nNJ2BKtajDSObMeelDR48TpUnsFK6gaa/TXQfuIkEgRNUh9ZtxbfL0bMnPUnnmo9fsLcJjUcqY
LGg+prNHUbXDh1QklVW4kNVbiLCW6rU3knh1GJOBHwgMkj9urV3uupum4q/maHJwA5ctyw0vOXOe
WT4Ito01vkWzKKpeSRI7/81B98eCdTnqLBoefUlCs0c5kxENrUUZZAmUFcEYkWs8UdtQsQ3MMzPR
/jugAJFkcHU470ZhpdF8XNeMYFfwwbmTX2SagnP66Ju6M8P3lApSfGvzjmXJlfM6C0gmpeHUXnJg
zg7Y4DlmQle5a90WbJmRVLA2wVF5RKGYWIzmOPzfly8gfvXbFuDK4R8mxYjXmTMwnzRXeEwhLwS3
Tqi5z2BmMIm9uWJjdERkODSlsL1IPGNYGZxHC3TQ5nWnDPj/DiRb9wk/gRgJo5VpYp/lRQKvCCvt
tB8ZQ8ERk/WnFdCk5RLXEzo3ZVPrbcX3mM7YxzdQ1IDWo+MGKFOVOke/IlmDBxFtUrvFp89cfPac
48apC4T8mEFdShNyMlsd+dO+cXUZyqnIq+NqeGG7NvBRgVIrs7+/nIkxu9Cs8A84zlRFH5tH4W3V
GrfYlC7kSZzEEWm74gNn9N0qZQB7z31vxxkYRdQka5Ul/NXdnhVxTdlsM5nT/AR3Oe+gcQKTVFbw
HUgRVsmZ7lk94tMpX7FlniNHUvOsWKAr34T0cdlcXmHUQxDlm4AJl6GbZwzZbqOYI7bynKcdbnzJ
GcdQZWwez5afr0RjBJPabj5jqF3KfwwD8ltgm5oll+WCBJFw9um9EK+0N7eq/40k++6jo2kr8IAA
3jREz/oiT59pqx0NQOQl6s2twA572BiJFe0GADk9JRMQlvoHVOt3A3nURKZzRDAjBtSiv7phfBQP
qkiRSX/GYhqRFHEV/f4rNB17BLUk+cRduLRytq+RSYZhDp0M+BgEhHthlXUWfzGgNuINV3iD6s2b
e8APpXBPC0fNPy3Lb9gGKyvNFGYP0TXW768no2MjmorQFEmfOzwWqhBP2FhttVrc1Rp5dvRHDA54
05HI0LWBhObqoZzja1w2cWiZKOUYb6h9To4kZ+shf08JHqerDGXK7W31EHjAPh6p4DHlhygUQ5CM
LpXgHBieFKQ4i7/jz6fn3oYwuP6UtKg/4AWNoF2I31KoR682JKxDfV4CO1e8zdjaHl4Hj6dFQFip
SLBWRTTlEYkVNYdkBK7qUd147YRudUZUBbXyayx8Ld2Gd3qlMqw4QzgcGr9JmR1apqdX959QZ1Co
lwyLPLP6EqMLexGyJy4khgBZsO4PH5SC2ro4iHuu5yAWa+glO5aSaO1bSGRx1uukhPCUvamRKEEP
HpLcCudE3nECEJN6EWQCX4ucvYIGTT3oLrwIH/8F/N9eA93gpMsgcjConHbBILcG2g6CiDG7ImBl
kQGidYS6QXlxGXY3AEPYw925cu/dYpQj4Vh+KN1zQGUzALB2ii+iODBWgeCjHPv11zFEw2X0PFkt
pbVg00zP8QCRvrvuhnUlPxelCXCifrduxgwa+mgFTA0MpcNTtKpzs0Q/rhMmcgBNfb5PYmc0GJZM
uxe/7V4Uf63xzlDD8PU1Ec/Gfkt+RxAMQeaDUUlx+n5Hxvg1HQ5MYt090Hirw0s0Wpe27pBcT7Cv
8BgngwV+OXu/fRebHRzg0xqtceGXDlfdn/oljbKueBbhwmzpeqleDSuGpi3xP9B7a8qo6kaM8xCg
Mne+KsnClpFzVMwLM3g0YQ2mZvvDdys8gVDvMIV+vLXeiMh3nUiBIQo99YCir3Dsxn4+j7eYtsxD
t4LUMwuIAnkNQVRQevoPHcAy5tQW3wIhRCKqMRf2Ru2KT3KAMFLzOIErkJJvZXQgNejJjBGNDtk/
lu8QVi8qXEliKj1u482W9EUltCiEZuFzlNgQ4qdACP4lBujTmG+st8PJdbizYFBdWoCvLNRbnMVd
z9S+36fI+Of409Jn/4CdWN8mjnviGkuWH/PTmi15Jk3/SNqm5yzWrGlaGroqbaK88f7dnRaP8myM
m6dBpk1NcdLe2NTXQO4kx1mOAru2IXi6knsm/2iQY9Joxvwe+MIVgci5KxQ0/H6IrF13viPYGKGG
x8kB6oIHYyD7sJ/RZhzVn+emyfsAFRVOIuZXo8+52dwPg+EZ/T6WD+5+X3xTJvTpZTYW0xzuJyQQ
GbhW1oq2eQ6Sdfs+mzANEJXQROmqPedfkRL2lJ1yxk9idOtWwvYgjac8slEelEP50yTTvhNGDFnE
21FCyneSNIkqi59aD2UN3pcWcszJvnG+uS1MLWR+v87rumjWyIi+r3CjWj9rtinhVrUCeXrTS8wV
4g1YAtkve+0jbIatK9uHlIp9GODZvalgpdRepT6pB2eYS6EFa9ZwpEVdymY6mJ0mN4aAP5DqyJI3
BHf8xU8IBj55Ivn8LtngGSlOcu4ZdtRttp70GSSQlU3X7x1RH8WQIs1CaJmlFqh7uaoo9zUMvvpf
HVA/nzP9onwMLBOzKgONFQvfnW1d/d0ihhuIv3/vsRNWsp8LtIdmFbRswcuoW1Ro2hIyHM9z3Uq3
83zzJ7J8HeiitW9s6w7dEkgXcLeW24x+JfBjeqW9zLAEbUCqMKOJM7Ema7YMuLbDCPNvtRLmhW+n
LaRvwVzSpqthpaQHwMuVNalUqNGPE5Y3npmjVGE4SVtSlaNxNkHqnvGbbLOpJzmczprMnvfo8LzK
z57Q6lLB64Sy9S2Aznkj5qILc6du9xOvBfcm+/8DPhPzued3mxFaj5T+AcIEyjQWDe9v8DsBpby/
GO8W5CvH3y/rCRSB9pIsWmZjuxNAH4+pN6tH9twKM8QsfovrcJzjFbSOotFlap/AJFlijvlufhct
oklOh3/kW+oR+kRINTyyqWqOj/a2NT+dzPOASc8uI9reDjlI5MzCt88Kt3Q25ESmy2YEfnwLy4r5
qr7WSgVSR+TdF0ZoA428h/3L/MILf9cPHy6t3fpSp8UOKflvOzgOY+t40lnMyURxbv5AKiB96cWQ
oP/LcfrpQh+amm35kNyfqnsFe6tj0AodQm63OiT4ij+J9VYNGxvSoS6/Lwxq8HSOvBNf1RNrH/fk
gF9D4XIlDLZ+CAoDr1GZd6S23gKIlu9+MD6GiWs5z2pwVsjFYlikrTGJujK0PY4hmCZhF6yEmPeP
82eoOPVabr1/PKCfSjRL2fvxTHDHNOZIdX9A7KAxjOVkRU5x8zEaySUej8tNOByOCG4qcDb6sXpf
oLmVlkFggXvu6eBCfHC+odmWc2syyqzGjaEUn2RSVLQEaiE0amR2YFMG3CdFJYYOgOwaVuxRnTSl
Mfz9MEZBIEYHJlIE/oOmMHgNP+J5xW+enH/VRZ6IT3GZ7GrL9I6GxGFnED0GEiSPvDXBm5U9ylR5
8/JaS1Fppkgyf/dggFwKi3qTUNxaBpSedyd0eNjtSsOOrZM9iZbIG0GG/aSJQykuhgV5ZOUxRI+X
GpTMKcW5vehrlkbHhTS171X+cg/5Za248fkOVmk9rqRntwiVLBCRU4QkLFnd0VZpx+OQf1/HZ6GO
JXnnBI0CnCSj0480R0PsNAo20rPKsfT1MoQHGyTaJ8hSPb0/2fHjv4TkFeUjYgpaBkBdXCmEHpN4
3cmhwWY25gpL2Ut4fxMeKDd3mYV6dnxQxsn4z/Saax5tNAhBNQPnn3O2/seNi0rUq0dExZiSTbEv
KiwTgijMOMRO2A0/x7ZylCb1rgn000EqwFPJ5bOMxBEt6YHOUtIfWs6VezsFPBtuBo8mPyoVdkWm
QKWhp3eZsM6YM/6HYK3M4EtSCP/HDw/0SV5oL/dP7W3nMmkXzWbZAYOgnXr83janvfGKp0dFKt+E
tZnNTbRczZDUWK97OJEgXAEhING13la7OopnLaUOPbJmI1Mw3XMSU0b3ODevVoRZhK7tL9l/sFhl
D0rr+QwKtvajBbx21aQaQg5oTru9tsYzzwWjhREJ4UApJqO5g9VA3KIbSdSlRy1oJWc0wzgBNeTk
zuR448oWx+3MnrSIjbmPlX6+iKeqzEsW38qSMhItLX4urB8p+iCUJQ7MGN8t0+lHR9F9gb/kbuiJ
8QAvxknhlylJ5Nm3QsJENzbT0AJDfFMTpWlUJb8pnnwdz8yqxBAZcXnS/GDDfk/VmAK4N0mIlfY7
4LHUPEpg/DmTi6DjvvFByLE8qa3YHfIMuv0gkCB/xMFCdzKOTvJiHMOUkpaZ3PiPl6KXnsdUBE5R
jF3RkoINBFMhUpCNvK8iDnMGKmOTkwnNsF5L/OrFlvcloaNWJf6adJE59p4NENiwUMFw5eyaNHyK
yq+K1fuFHfynNGJ1q2H4DNN/wFz8M//T/PjoMlXn6VdxwXR3A2KjU9Hg2RKcfECFn6fh6WCKmhfK
oxMTk0tOSBuRtfRm9Ns/dFnGYPGzUoG/e1nkrh8/PbOAYHYj847jVghNkpsVWmx8PLSTEoywlR4V
8jrema/R9jWYJzNAfSwZ4QzZ1yqbpMRGy6K+jcELbmTDDbx7tTJBn5h2AaO+9PAXEprBwb53/MdX
EyH4Qhi3rouoJQhswfqWodg+c1R+r2NMF3mRjbOXDNWUTfRx+EQgSaTfuXCIr3kdKDpmRwmaQmzn
rXXXSVMnyHEPPaIGQYN2NSssYsq12knecq1vWPBAiXhi66W7L6pg+W6AODhmeQTUZgmaGRszs0eq
rYIWDtcJ1vYlleJjWVeAhqQ8/BeMTpvlktgimurvFqpkPJuvm86/ofcbcIApnImfDj0HnzMtuPzS
QmVLpU+dcfJlyxqqNbsxWICJ1ElxNBroudXm6qGetdd1JquZhMPRZ2c7C8Tm71e0LRqEZtQENiHp
18gwx0Fp+ftct0EWz5UiVBAarP79YLQOVbx3ctSvRVZtETpk3BY7rO4RwpT6aMoZCta84oxYKWRG
cqAtkONj6Z0gxZkYIhGDBTTDlOYZzpFQTt/6kiPEzK7bbxwQibenh5hsb0lk7Dh3V10xlVT9y6b5
l1Rt8GgRMtRBN0E0QcIyDl00YZCI4cBfeWv8gtjACfBjCX/rn5yGEDHLrMjUpjWLSz0OEbev1C8b
aYzoLTagRu49gbMxpwXl4ovnCyz8A5CslLDzm70+cur5ISYdyCQDoKcSGfGhf/MP8guLJ1x6cYDV
d5xsHtJpf2A4Y6hbsx96TjkDGWo5AnYxUHuMQV3RRpIhRACdJ+2dCDnHgWn2xabDKF17078Tgg9N
++DOg2JNbjZFHfWCYSml5qvCK/hOsIJMAZ2rbPeep43f2Rk2l+NenuqhsfUGX66UU49JIOTMvGEP
F8dqQoZ04UtjmhnpdFDZ8cDknZIa5TJPVdHTCHuO0+IVm3IgcavKqxuiEnfrHfLz4b9PXBt7DAPQ
bHXzZcB1L7ZBVBVdJaYF2a12EqUa/RrCPIrEc4LBK8etPlVD7zd98WcdkiM/WZwe3FXYKcAzfzsi
1V/HFmNwCV1UL+3kX0EKtEzdgQtvcRoew7tV92GWDr7+6ib6B/mhg9EMs1eecomEQKZcLv7KSkC/
12fVv8y7giag+peWglRuymkhPvM69p11k3r4dMfz7bYuC3mBSKzpfMpLxAoKns8nyrtuluk6Meet
BHMsmosV6BYlBDP/akkmLeswX0yjhdck0eVzEIYGbAbgO1TbzhZxDO9vknYHBObvR7X9UvIbr2Bp
u2/sUNbzEOexICJ/cNfxJ8W+caLzxDpERB62qd9s+xunfGl4Jyau7LKEZ5vznqn4LNEyEoVU4Duj
eNlg15bVMrVpvvs24ky+X3QmIEtMyj1XkA2f5u3B+XvgDZU7eGkZZDIEuxHWgenpa31edpDVHECk
QiBQqu1iuKaIdMlwPKmxDhLDMum2s59T1OHmLYFYDWLIVdmqEx6L3JtWq50jBPnbt8wK8G2so75E
88yiBmtifjrhUSbAI0A8Kyw8MGdJ+jBJzypvIOi2YgvD+MSIZYlr4EozjlkPfR8Us52MvrPbBbSK
9TYV7U9phHnvkXgln85pwoXMHeXFt7GzOKDWSV5RadCjka7ITifDwCRjkyJ9sg2Yz1COGwWSo1Mo
Hak5VlUz6w3KsRVmtL9lRHXCra/XOFUcjRjPXiBZ48z2slgz3v1OoDZ9bNdMSuv4JUqWe5jMHQCX
fGGf/AqCtt1vYygJ6TG87FufJYNza3LorfcB7UyU67nHI3xACa2IOsYzM70Msdzkrc2ODvPubwO1
WRlKmq4ZWwHS64150WklBUWuxgYFzMpuFXNX+oNU/ALVDFKbOkHFyuslC71A3voFYi7tLmDyiZFK
kbCEBXsyN+hdh14HT6d3rMbL5uDFG6MlVNlSeeAkFFS52CX9K0fA0S0PyZ1YECSjuBV/WDuWG86j
67yHBXegRYnfMGArvb3xScn8UeA1AV4of09xvotD4tVNIS55oeCXUerPrnJ5CMZ+Ox1T4G7hjt2o
hvrH8vtGOwky/F/jIhDh9l5putYZqtLgXV1POJjbofpkBk5ivGUTNLakUAa2NE3DTRP8h8Eg44bg
swyoLpl87PVaFLIDE+XHASE7g8YI5JiyefLe+MV94TR/vwR6yap5WFHLdL5Gpox9kzhTTKoAOBSY
kT4KnzGFRccwc35f0resOOWrkkZIJJ6jvndpsTLXGBaHOYuL9qNE8h6Ef4mhEz4A70/7lEOlhhHN
k4ND7wT+R0N/fN2CBpZ3cTOfUet6sLLwLmuRZy2nNyt6LQbE/vyUwY0gU7VH7wXT/lex3qCcreS+
5vdlwWmz7sRP7+TtXwjRlf/JNHpHl0NgD4IYbqcV0wywPFlM8kbRBju4wtIWnL7SVS0iFXHXM+wQ
KtdjkIn+4qPIh1UYA1rGyM9X/eZHknRYqHsWHyOLi7PkTa59pIuw8N5eediq7OYKgito8+oaNifK
hW/7VLf4dpMFi1y0g8ZIwsz1KQnGaJGRkia9L+v3GzWQuge9/BudmuIVhYd3W6SQqBO5pgK6hn0X
GpYYiAjUaLCbjXXa00rTmE+/5BmH2TAECj5BryXB3r7bUhFrGOl+41VYDmb/WChXuLR4Sp7sg713
7P/Txu9tK7GBeOHpTT73P0oRy/mYNZP+xjlNPDPPEU71m3twjwIfNZHcCbpfInQHYWTPA0gpDvU0
gy2rCatH8ZxKlmyQVCtNs/KXHSTqKOwa7548mWGZKyx7hKiEB47DpVTqZFarT7uZH+8UV2Y0Irm6
0kG9J2fhKa9KQjQlmS/BGOnJTOj5sHzzgAFwqAsp9haw8BHJl8VL2Z2w08xAGhXSztN/MlLGQxx6
mzFyTkFSSdvulRSJvHuKd63LwRro6lJJBh7ptsK/GAlzlaJwzvNH8cSeYl4ne3g4XfVCa7l9IYKF
x3IFKW/sJN8v3sNcY32sf3ZBM3Vf9mjbLZ8eqCdziOz9ReKlv/JoCpWD8xDa/ZI1zRJ3vyOGFtuA
hKgYHKoS2fxv0blMwxTx1BKkra1+M+kgU2p0yD1HlT4XXvmWsmwj4nXCSSWm5RyiedT11KV6R9OO
pLG0iTd1Z8P2pExwr4fDmJP9ygB7lBNlHoQ+LrXUrHJxblkGhbZbdma5w5HE6V11LRXnzqOUpzJs
GGDvm9aU1xVxg9lhP2arvGavL4yNtg7vxw/SEtqTWzmvShdntw5Z6QWQNBcpIVaCm/LfH0JJoRr7
XqfZxj72COap2tGRI24vuxEk/IYTFmiqcQNANApMQxzP+UdvmHwxJn+CbtqF4hKelejgLFXZZ22N
X1JRhM3XsIZ9qHhTvm6Rv9PbtNwVfaTbZIUkiRXAl+12SYlYCd+GbT9Ft6lpghJ5xVkihmWi9d5n
Qi5qXisosx17dVFYcbyTupDMgnmvB+PJYnWJbMZjn13fjyykQwsd9dSakSu7zpTuSMqxgvSXSEAK
5jGgHDxmeItHr/0iMN3wdmgjxR9l2NdRwBegs6rJIkEccxoyC292zK2fRhY/i3iPMaZZGFv9ZqtC
tk8u4bS2EMhRsBEcSXrDJCGZkEUoZYq7tjsMvNdbZPVYf1Tka6HkYGeLULOa+v5MNZgYWlrYmCA1
wDOL3pZbtLH1amUicUs06tiQwcRIdY59fBypXrvLNFMM9k7CGewlKv5CoBlDSrm2O/IWoLtNevez
+akhXqCWYRqPKtVXz1AVCWMMehnbeythhgyh1dDv51RfldTGWWYHWxjXpVxdbpVYvRJ5Ce9IJAu4
mwH1jiT5Rp2uCxTxB+0GSTJz8xXDtLcP2EIGAp8dZ7JvWefqti2uGq6KnRUPPBBUJC9CpAhbhQGL
oLNgi2vVIABIiJCb2TdoMXwnAC/EghCmp6ROCH3o5Co8K0bjkRC2aK9cQUgIaib/gfG5YGE7NzjA
DS+jXCorquTFidfz7Om0K6UOJb6AbZ0lJkKRhayV5W77bwyszsJb8tw+8LftQzNSH9rH1JcD58Zx
0Nya4fJja9LE3q3VRsUi9mFANvGpcfshBAFW+6UxQ+x/KOUl3OOLF8NyMXAo/M8f2/hEfOgWLw7F
9kLJrsbmDONCBbVvFhRsX4deZQM84O4E63A/0O09h6dTbCXUoG6f8RGtAZJPT8hY57bkXJy1vzBP
ukagOhZkIpaaEcUSd2JJbLSRryi1lvOFix6VAuVD3rU2uzxv6bFH1OOPw44DuGvus6Fcyki4WzPr
zbqEfNKtg+Pt+QQnFWJra2CLZ9AFU/cYDDflw/0TXDn3H+D/qiPMzap9KNek5MK/mkmkW6HjGbzQ
XJNxogMMUgOwRJkirvBNHDTb4Z9meSW8JSoMyg8NsT5c1j+0YT751/++Tt8Rtq3VlrjYrO3ReDj7
Coqn9JJ1nrrTSPzlKKHUGH4pj6C5dvNjhYomLEfSlP7aZ4duHxcblQ61jzx2rwdzsXRWb1Uxf85Y
r5RgODZjTQIoukVODJP1eGo5vmb8CKt8WrDNDK0j7iGiolEoQHiT5I02GBmmoLZSap5WdAuKlV8P
cThLxN57ETHQg3iNd0pdNNrQ/4bndmA3O97Acn84LmLbT0Khkqgugw1+tOYv7vDvw9Sq6yA/71tX
I2LOgW8vWnc9orXE/4HBMNpGINKLO4e4uOpTX7MkaUjkZ8HrfK986x0hHCo2oMQtbBZzDZG/zIT2
GHs48NQjTXy6sjzOGE1ZBtT2Nlw05xFFx3g/VjKZWP8P/uMP5ia2o27wsoSGI9O/VY2RBDwFId6Z
/yefC+9+5uHmJR404D8ePMAebGgIvz6YFmxISyX9Ti80R8GS3304AeP7csRV9Pj0KOy55HukfYaZ
Bow4N9EnpDmJykchnsMsFjQ+e1NaIxmO8lKgTe1uorcvWf6vNifz2sdVOPwKfoQQ6u418jVJuj4f
XPI5pcEY0L/XVmnGgZNZuDOKjxyML8MZpz1KLm9F8Sh5UNdWRPQ39kpytpWhdyrapXmpDzQY+LBj
ySU6nY77ZFVwxFIBbTnAMbY0NfyeF3t7n7UC590lliYyid9k+rUNOu3lM0bBn3LZcyxCyeTPK1jp
J89DgBdjJhgcZ211BhHWu9n+pDmr+H/g9TgKPhh3nYpKm7dETuUc+0Z2k4AhLEnv+ttd0B9v9G39
GoHl5xJnJ45/sVyinmxHlg2EaHgL3n4gxGtPKEUZrMGTbBmGq2yc7f/Ocb0tBrYWAJrMm5Q0WEFa
LM4WaMIv/LxzASZ7FJOP+cuYjOLMx4gBqjVNOnPBRlLcJ4YJ9xUnUXL1/LAdAtcct9t535rgqn3K
KjELYONKKyOW6C2etzLPR5035cc8DhBedfwvSm1wvlAylfEfr5YYNOwE0lFHY6PuXxH2rEn/iQzn
SRblfTwXrYZZUF/SAU3cH/BvKaaXz5S5oOsv9asEZaUy4/n1jbmWNopxwhVPO5kZDjjRxAJ9HHUZ
r9he2NrtftosHBe5McSus0Gic4ODclpIrn2rA/Wg8h1lS+lAAw/yjc7ipasiQuaTIbrI05oe34DU
N4L+DWfhNSoLR9YR9iGL3ynOEJzwtwU13CVcns8w1wB6qPo8dePTXG3QmfPddxXa/m4ciZ/W3UVF
ASOrrICzCDkIr7Lxg2gpfH2g0fwmZAJ/acchOdEgAjQODPC4RNnotfBpio1ti2+HnPEQP1pcXaDl
6KIAbpktYVjcUrCABAGjSqId123Kzgkj/2etG3+K6FJKgkzf9rFkQolvnWQA+9pi2GcHyvyqUxLL
XFxkomu9gLlGv/f1qA7z3T5DOojG7jxjWc31BiaS6YGGMtjhkFQE2F4P7/vlk9YQJJ6hCudoaEPO
2RHQVDd4GAPKy/CO/S6J11qap0ijVJt8+vw/RvbxrfqFOiPCgZUsZ+ye0cjYfRL0N6Qp/ORL7UW/
dlSXjGpdOFE/JMmCXfKJwvEHPDiBiTIYTaX2qKWPdM7BtGCmFA5yLEcy2FNszp7xPfvVGfbcyN3e
r5ZwJk3/hC1yf/Suv6nuRgtEhBnKyhtnLsIMzCe1QogrgG7vW0o4xHi3jTg69vN3vCUUBve3+T3z
m0jR3ez5G6PYHV4K/P0IlMqykgUyuaE9bkLGRVZn55ynjxXYwDOMSmpw6rrjpODENcK4ItZs60Ya
3A+Fpz+OptUaDIkKW19WTEjiy5GCq6xfl5uM9QLGK6kSKaBtLfRKzG5ebQA=
`protect end_protected
