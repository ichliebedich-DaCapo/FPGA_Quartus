-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Eed0g+1bU/i3vkBOApnjTQJXgS6Sy9KaXdcBLQyo/BCRm16sGwQRlRGtI+3sleu0wsGkFeJKGPOv
csfiY5fIAsi7jN3HsYi6aEaTmPaalbo/XOtnnjDQllVmlxMGmgikhOuuBQVwJcnLznu1bGz8Quh0
28XVrYDKQuCet/Zz2GktS8Q5PFsKLvwEHSmpmXNYkJqPs30H3v5KJzIcfTpQvOi8QrbbQZ/v1ODi
uBk7UAc4fmFXUlaW2ywEXZbg3zZ9XaVfVbhyfopQD/clgqHQMc6/nnqGZM3OmjI2ZQ78Swd9roxz
sq5C8nLncJvFM0yB1gIrB9np8ggrbR/DWuZvcg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9552)
`protect data_block
7Owc6yrpeHO1yEslGutQtwLANcWXmRAPNHr0lPNUtEtqS6QdKzpuho4oMcwq446sFmxLQ92XwnDX
xlc0RZJXmWgDb34ARWOplhoS0uCEWdmYNgMqUSXD45uJorAVSLmIXTkXTQpyjlnYg5KEuUTxolZy
hEun4jNaTJtfBRdsT+EqtQ3xBwcMXcx4AvR1y2WCYoR/FQNhpO0dcR314+TugfOJMcx9o+JQjYdP
tOpKslkikT9+IbgPexMVdMFN2jZY4WBy5j8wtFsiBBH6cUIhLvCXe4yergd6j6rQx92qysFfwrum
NknYPLjXRhEBszB5rvuXXK+tk0vv+0QYLlFce08suswiUEORIaNzFzaueD4GEw2CwovQWUuDmoAF
vOJD4mBT2RYE5R09FkfUCOtsqny3dxH9ijDBMN54YmP3jLinpY5L2ti06RaL8LMl5fK7VWDz+uzR
dFLAe46UJihT99KsVeMv6n97KlvSzE6ECRIXgLEhmOL1Xug23itduJD6wyqKypF3EiYDHf9gugwe
tn5pkrsqjH7zEvjc8yX/HvXq+t640F1J+YRknAQvUsnPXtlrXQAYsYd0FH6ZqD+M2KLBjUAd7QpV
E+VcygFCTpgshxXUgmmiV26WZ2pIMGPs+0IWbKLCEQv7/vc8x8aJgqmlMr1jRJ/tTfIGDUa+LILI
J01//+xH82DWqx4DHa4qiVYHrC9qUM608SFmTHn2GYS19weDlzVba+2q3iKHljfqQpZv+1aYaPBj
CaMjQazLml+0UkUb+7o2WDUNcO3iDNCeVLpMBRGrTvXJx19XWZm7vlKjS/ekSPDcU4cqQHkmVN2W
FDdOd9Ll7+pVucJG3jJ/TDSZu13VdbSLnQsqLRLBE2Z9lLXvsmqalHYVYSe8Zl86ouPk2PkfTXwk
6vaSWM+q7ZEj2Xo84nIkfk808A9WIn1I/MnjRQ59ouW9b4LtGw6iyUfl4lsLwXoCfl1dVlhGtdgL
Avfzlr6MebRk/9ZvgFPEjveZBST1M75WMq/r9577vmnAqFq6JEXAwhj0v/GQqWfzMCSfaUiR/2z6
eEjkbR/Pn8sk7Evt1M2Q28b5x8Q0JzpY+GE82cn1mRlEDn6FAs0e+9toNu3troi4CCot48ejxs74
3bKBF8YIWLzD5ORJmySkQExu5w2VOblhTlVbBY/puLkSTGJvJ6o2OV3vl0rhQGfxL+30FhFoj9YV
IjJmUvV/7dor8gJ3qNb3CYhIqMHfyPNLMchzrYqK5EF+SLG4Xmt48BVbh8fOgLcQHgo78B3BoQMH
qS17eVt5DHGeXdLiB5U3hsOUgOXbz9M1nRv1mNa1hx4sF2shC750pV3bGcUFMbUG7aoMKPbODiRd
UO88ogd90PqhMfIn90SiwCUzvkWbm3ULA1rKPbFZxFcTEzPr/x5iO4qZYWDfluZajRzL4v+QKhEc
1tcfonT7himaTZJ5fEuAeOm7kucizS603RVrkRLPDm2056iuXUcyCt3BXB5eRtvwAkL5/Yh+d2KV
/FZOHTJpWv/2QWAGd2sylTQNEoAF84Dksoqx/lZlUO+lJbAOoMLKX+XJv29WV7crjiPtWz31hpWa
YEZK+vTmvyikvWE7jc0pD5idqiY9j7jpP+S1+B77wX4+X/NxSDhxQ6SvI8Imqi613Ada63Noz/2p
HKbB2iPvwkcTsJfzIl9PBTC0sZ+kceE10xN8Vsx5e+hiwkZX+U4LAJNhDkMNpGzsrTvCM9SUA4R5
qraS16NTL1qBfvkPWkGXbKURvi2TVyXvfTZtqfg2MDFzEWwyY3+G+6Qo8P17vwqSpriDGLRafOA+
GarztM6uzgMR9eYjGrphv6+XwOaH6aoATwqioLG5yoWgzhIJ4U4osKmgL8aYDOxdUg06wOla5ZW7
yTowo3fo4A3SdMn8B8+FEgH5//m/wVdPtzUov6oAY6WI8OFmRk5hFh/uDbEgzMmNKZBbQtuXh+h6
+uW44bWesX60veEVk2fGJGwFViwdNrMLsu8KrpHpgK0Tve/H4BEJOiCrEwd/E8duiaYOSIlbrtB9
2ds0UF+tsMh5Pk5zo1jMrC5kuME6PN14HVuMQQIVU1JyIbpyvyOjS/nTcJUE1T/Hw0Wpdqk41wFy
g7bSdwngpnYPTKZoC0QOQLYIYInW+/vq/GCEp/zdUXmwsaYbI5L5oiwF44GfHa3VpUXA70fQkqld
QPOIYaMTiBfOBjhrM3M3rAXQQq0wCpmnZ2vjt2CR0YMzd8lpK+vyNpHaLTRhs6bbzTjg1tdHaEkU
SN9bO/LTwQYk86I73lSVNW1w3kFtFXqSYaHMOrxh8tPxCxte3swjJAJO2YxDzYQFPByW+z5iJwsy
c+NyYw57TgOMneXHJjqZscue1WrH/qW9qkTWoWgeQXuGNLuBjhtYImV2BHvQPadLrF4ead4wAtKF
SS32e1SPik1UNT0y9JvckrciXwkQv+b08GvIvtgAT25xABEV4z/s+6kEzy6ZQUgxlKMsA4WYJBiT
FiQvLhrOskTrVP5LE8FIOOcKR4cpqcosVyNs+ed+ND/oCH5MZBqU+pwQaJehduZxFY/47AcNLpI3
sUr3PKn6QftFQKKpyeW9N6e+PQwyQvYcMl1Vtd0iJKrmHUCh81gSZ1oC0TofdYy/eB4odAdxYJlv
7xAq6cCvQmTmag7EO4qMu6UYK3rJLn7bKMrAMM0HEwb2qe+zzrl+PPILGe7rZ6EshVZv2opu7Y/5
Pye4PSckU2/t/a5gzgY1M8V1I8SLakWbAbhd6pTAjUSW+hUAc0IotB4ITwfN4VgupkZfk06CTfHO
52MRXIpOTrOSYgRMWb+zOTFOiAilg8DBmjbQRB7OSnOrdKA9fkQ/snX1FUay1KA51Jp6hyieJgtd
k5hLEj8zfmClg06M6NakwyDacnVoQKzgs8b5os3C4BFfMqvqf1VfDNRna4S22hJ3giyctvZi0O/g
D1KwA+5nutxxjSEGiKu+m/TfHTTxxmonys1saME+4clSRN46qwaDhTL0CFVwQfsZTI+6l1Z3wZ/l
DBwJnqIscqx+ZIPw3JrxM0n4jrMCfns3qx7NjntU7b8GRczN644Kz2JFosvim/dhpj4rfzLKfCij
Fh/HKKALmq4HIkjZNtW2vNDIsbYv8YHR3c5e+1JtIVevIRKPd8xfdP+Rp++EX3VtM9qL3PE0VCS2
py43gLnldqrszwBSilXreus2sRY0i60C62X24W2mIqK6a8nXemiK9AjzSohHA9vDuLFrFeVm32ln
+2dofX5WXlTkBLWQZAsCGjPpWmUfayRxYlJKkbi+gN5owe6uYa8wo+Wwng8JY3a0vFG30+bH+q5s
WfY3F4SA5+IEeYeS+tR4ekzjAloipcuC0+t+HW0Za0495FQ5XlhD58/rY3mntgC1AzX94NCjUUOV
Um67/DsAPtGT5/X2hoEzhKEBjv/YiZIET56IJZvh39FQlWIILUbZZMxED1jddPibCBR/WiSZhQ2T
3hB/X05F+VtVTu4+sRubPNBD8axepFVgYo9P7UFGGhooknVF6tsJOJOLrBene9pFuk4rfn5YW2y0
942AsxDkcYNPlJmyMtQB2aYFWfgqp98ZazgFdXzGiy2zn8T1VqNkI7/fCm3IUw3KoKrY8zW5Xrs+
+6dfcyb5/aZPXZbtwnKLdcy2pdgTawUijQCVaosoPlcevdoO0nImg8yv7yL/mqiWDcl0v4u2DbQm
zQzs1qW+EROwukCDMFW3HTwT/fJTdf8gLH02SC7KMHHAXXYz7xZQbCXbRYw468dgfgjek70gCqHv
NHLKsjWw71sczlsEbzBhh4tmiOFcqZmsZusAIY62fWMkNK6W35cbbERHZYQxYag7Cep0DRrEAJ+Z
qccmtsXB5DSeVryq3CUJChrozPH7+3+i4wz58Oo6+GLkeTxgNhVH0dtfaXxPVnEHRUFeK0QNLurE
64Wkxvd4dU8CzbrokW9+HNG4EBWtnMMhTr3V9CPPH/nYCteXSVj6eCBY5NZ4EbNgcl1W765OqdGE
LARN/VzcPD77ZonQxRp2/wj4QTBa5n+349qtrziCZ8G25dVFVTllNE+SUvmzaISQ47oX9Rkgx0wS
/hque+lyVl5cSCdh35kU3GsD5ZO7ladHzIUK6hYBAmK0HfLHT16UU/X3sHIVTkGaY8W+HqRvbp9v
QJ6YJ8d6AdLEBE2M8iFPINrqzQBb3Wv6bvGmpUQPGj2jb+PmZtWbKoy9ZlEP3wqDbldppMCFYfR4
MzA4A2Pu0fHH8x0LZGyYkIflm9I00AgrePXPhwYvDCyOBTsbxiZfpLFv/fZ7QRpDHfmnuIiVy7Ep
UJyWYnX8FgL62qIQTLd49EHW0okXNsCzFC0xs9DAZIMh6rjLhStfQx3/TTtbWxzl/FcTxUWFUYK/
k+5oj0SzY4t+JOOOY7z6joD76JMJVSoHo++BtKvN6utlbA3kDx41UVM7Gyd/Lz9Zitp/YLcluz7Q
kkBgOtT33UsViBwNR5HvlE5H81gsTi/8i9+0qDDKSj7u3Sc6TXZt4VgyxvRRrZlswEN9OqWHD1R0
/3Iiik39BUzumDAm1MwUWZxDSmM9MbJfjNFTyyFEyZiTlCWh9E71iyyPGT7SbjReAUmxUPH84aMA
3krHpv5m1JfTY8vShvgZHFP9VCnd9zrD0M+nxuce33ZGEnn0wWJDXPb62v/3M9VMXuYvbU0DDPF8
TQ+9Ya66/j0+cbvBaQKJ8yNnEf6xAPcMqwEJgI7JIZyh/0IufXzypXxURsUyt0o0CQSJ8AxQ+FhK
dXBs0rxJqgRAT4U6LyCI9j69ECjxms0Cu7S7z1eFaqBIR947DXoSgKyE6vbUBQGbrBOKQybR9Bj0
/ilIQDxKbD76lzdtVr6bQNSG4GVJUbsqyCjV/V9mvAEI6iM8Kx4srV1L5/rIONXe0DpaANczOGVc
Q9HabjA/QkzAbgSxuNsNhWUCZOzXjNx/NmJfpDP6DvnkwuzD3BI4Y5HNiyyk22CZVvViCAHkbiBG
2bV5CHgDVgIR7Ty1gMs+RQA9A9lUebVMxMpzqMMaDsCbUqrILjXn34BtbCuHeltNIgkvW1gOvMEd
6F2s3cDPUJ2btA9hKs6P0Mhv5AW4V8MtUwnW8LGlsjzXSbWTJ63oUHDjPHrxM/gEKnxSgy5nq8de
wjWwNHafAHM/z/HdUnLviJj68OM227ihG3+bCccwG/uu/YY7S0x/a10nXTlDM2kKE+STKYGivo76
1EyYMx/GjwnbnpOCnAqV4FmMUtozpmWZOMFBee6PBjBJrL29eMcq7ncq2A7egbp5gbJaNVHoKBDd
81J8ir/Q0Z1dwgalkm0uHoJP8fIADT8whMjc1ILc3XMaMKZR8rgHQ35INZGrCSb035g98fP7M8fx
u3X6li4wHnTwjjh4srhIJaigz09svlRbNi/8jQzgiRjFpRI49vKx9m27tgMq7LBeN3WYmNnuJ2B9
Hg1FM6NF43qNRTJUe5UfsW5Lm9g9C6PlQBr0LZwJlTyY2Ri0O3QLYE3hksIB/7m4kOMZY+kJ1lTb
vZ/WO0MTuqBIneWYz8dnY/RqZW57sOrGAcyk7pOLspjHv2eNXT/Bxmh+/AYvY/n9N+WlGZ+XJKZ5
f3GT/6QcI73Dl+mgKsoUmK7C4RpIkhDE05Ozj/FXUId6AdgIIBPPNVpYyM8oVI6Wou9iOJOHOm7o
DbGAsd2YNXEKuY6z9fB1y+p1tCU8TOWWcV9cl8JMFfxYa57qpuBh8UQd+T1LP93RMk8ohDP5Pr8A
x4hP59PZ4Ye6Prsb2Yh/LkRYLsx+hjyqTmsX5b6HIcE3j1JseBGgZsuLNu3+hPHXKMraHyL7IeAa
iuoxpX7817h/8YbT009hkDSy9Grz3Nr7cvZ4hNdXj6kWF/BNsm5e+k0W4MX774Z0IPxyMreDwpdn
eahZTZ5lP/TUws/+gptFMqH96DtNVJqvnbcovDM0u3D0PMuBKi4rOXdknq6gDHayX/4Evc5fX0fy
9sS7uDfArw9rW6LiPksdYFiky22hjZzCaQEaZ5wngYgranGfO4rKP2mWHhIVLfpkKMvinEGDmild
B7n090Pu3HKuWTCuZeAN1nHjetnojJRnaUWNc0CxCYve0M8oMkCo5L7+YKI/cTVK17rR/KQQhhPF
droS/N5ilTZiJWwTvak/3MuMYri3KLLqKlnWQXnntTcALUKJdMLc9GQaOynIpsxHQsUUGw2rcxXF
x8l9MZQB/6GG6F3QxJfuxV70bNGUcCVQkX6QWSkVU7yHDnw5lbGFvga9UCEpxA4lJBHcPmHs8ldz
pBkQxDQ9NI+blxaYbreEI/vSSv2gLHdqtmJVScwO8C8EboSySLYYQelsctaTeD5lYbTp0xs5O/ua
1InosTjoKpVNvJdY4oEEKlf+08BWhb6O9YyIUmd3kbFRkkBVMVSnqxDyop8Bbps38SFZ6JU0wx09
eHxt5VxBkue33UKc1PIrwVZ+Kay8GAgP0wFoD/7fPM2t4iFWwo574wW2W5zzh17vO6qebEN8zXvk
uYdU5SGtGR8rYWbpt/iLq+2TEjNYRhrZ7fVfPZfPyAE9k6TuldjVDd3hFgDlBd5DlbUWG6dxyDgi
PEobsgt7VRNlffD5j1a36zEFSXDjMcmcAVljuScYWUBHa4rQ/fHjyYVjPmB68qA/DDc87jvf8onk
iWXYRxyo5CRvG8/q1ioK23aTK+9eeAQ1ym7poNaSJ9iIibAdAgRqkZkPm9YqWGmRTGtYr+0cDfcx
x9VjWHG9LnY60Ql1HnESNRaY2y/xlkdc5GhA/j4ssCGBfKDY06VZhFDsTYklk1BpMRfiGrbQ+lxC
nB29qH82Qtf1/IShdGBZE4ZYOBx97XP+gtxNLaAdOKg8EjuR74GWe84tz61NVQQpQTr4X2eCZ+kG
nLFW2Rmi28FwPcUlj2oHO1M4RtiYNDoffHg2wwWjZF8g7NvG8qYYUD63xB9pIiyMQBTWdFIpO7qD
jnEfrDJeEF9UrteX7lj7yTa5j+71/Xf0qIqhEiKKhjW1bUwAMy4xP4QAW7MYRclEIH+dXsGPKj6L
A7hSdJsspKd4mRJOedc15RoVYnlduQACj5cB4Ch/lWKw4bvt0inZZQ7BrLTlBFavKALg69gTz8w2
iT+O5Tq0/aHoSeLALcr/XBc6z7SW1L0tGJJtpaRp9xs9izgkg8XS3Aa9xj84+VJO05iuXcmcMzyo
B/+X2jGPVyL0NdjOTBD0nD68gf0z9xgo5KgGb2wIkbAKYct9PmU+mgDdu9G/C4ZcOEjSk48vlmmD
/qKaVnQMQNuu8QLGCMmVnr/heluph+tMI0nOzmJZAE1XqO0D6BPHbRKvG9er8soPd3zz3Aj567WB
MxD+rQ0qkaWHl3wAavp21s/oQMSjAXvswobQmw58H9N4Iy1OfUuM/fIhpK4hBQtn8jCPWIMWJ3Ev
o3mYhRG9gteNpG/eFKHVXSWoCazlU1EsXWKfYEO71Q94FfZocV3ofCYutHaDhdWlsh3UbIc3Olgd
aZi/JbzEyTbbbkvh8lNidu5T06zkc9QPail05RbDP5874G7XIRV4O3UQe5psjqvbWDbOW4xnSs9L
u8qb0SUs4tOLgp8f4rZCowRL9ftIdImsf0Dmui+CFiY8UsNOKrDk9PQfGuIoGyMSrMZnMuCCAoSs
t7m+2taw6DPz8G1oa2V14px2tyDbkraNWSZgwcI4vOgz8ByZLBBYTTbna4587VZ3wupR5/JAn4PY
diTtxRfMSE/cTpadlTMbE2lViFO6hdYYdrJTcdw2jOtRTmzvU4S2/r48PW3XrjYYO2jjaBnuIlQr
OiZEk2XG2uhoJRnqhTMXBejA0VYZiSUKUd4JqLIVYAC3EPNoMRnugZvmTHvtyL4kn99JJP1z0Xgf
QcuKmBLE24ynoaGf+VmEwYFMfRQPv8PiM6ZR+vXfkRegzm1JkYv4W/L9MulAdr7grNcD/e8HjbJo
nmj0QIXeV8dV12vOXJOjP8KbGPLFqabnDnOR42coliffiBDXUpXr2I1HNYZaKXyzO3hV5Cw3BNSy
X87mF2YtmksOkIH99IcyGrFlDztaQTbTS5GZKwXhrzM6OHD/nrRGZ6LuX6Oi2e3eeqLMteK1419D
1uDbiXncxmRqB6bA6Krq3BVcDoLn07t/3JjyNroya90ua70wkhfG3ZF8haPjiSD71sZvM7DJMG7a
vQn2LXIsDW5KtIgDncAZq8lWOAhzjhS39lcoc81cg9YWzqRXPNM3H8cid3Rmxqi7ZDv5PYfT6Y4+
tIkAAtnMPj0aRSufjurft4w84KCYvarVJo3TxplubbMrJcGBQkgvK238mZ82HtKs34l/WnlTNIKE
sugLli4FmxnOmkV7tSja6XqAoAXgCN3RSHmL0dSGyjB4CHGyHsUN9F7mqIP4ldbuy93jADFGERe4
u5YN3/0V1URZFuuWMqfT2fP2/sQ9SJQq3MsGqqf6zvUnrjoHKLDAcfa2/qmv/Njlb67qLyMgHENq
wlHFqbTqzzJFS1Z5teODewgPNIj8OWgOOw9gwYvotfozrIYPrgCrRbM9AyyWYZHdc1b2960fQIho
rRHnyjx58A6pYLQ95nAAkAA2HuXNJsZDWZ5lvtE8xKnkMq+DRRdbm1e1PN5gcxnc54YVM5/zCZIP
gYa3nsj49BfECG4Idl5kRbFLu0syB8YI+YsySwV3VZTRlxahltVoOv4LqALzdu2bvopb7hWJTlP1
Jpx0ghk8ZkycpMctMk/+330IXoywZj06W5cohGu6SW16cwIwe69kBB1ndptHHpISpkmHN0PIYdfZ
231PvjUdjZ8cpmFZcnRxGPM41mAlZB2ziQn/+iufbGNsgn8fXS7gPQYt+jfMfh9jf5UXicPom+Gk
rcKM3xphdPbXGOC95vnw3w8LSgrJCSf6tqCi1a0zcahSr4sMfcYXRp877w3x4iX0z7ZtZvuQSlLY
ittKhf+C65cJ9vK3sxKsAD1h3TCp4QzlJojFsoPYvJHplRsf8YTXPrP1Pluue8lpUTi3FVk1gMj7
M56NPPZEEvOL66wmuqUUPx6zIlU+rKxJHw422Af7mBsTYmvt4U9hUACtV8KG7R786XzHOkZuAvDl
dzib8TWdBiOMbnPo4CeY5gbpeSXL+QOYBLwfn6/DkKUJiCgQ4V9Ev5o6dkpiZVSG1cmudYNXiFAZ
Eir8HZLxTSErWF4cFS+NL8tk+PIpJkWplV4TPDJfq0n8ks46Re1O3RIc7FqRlAED7obfXPZG89HZ
TNMWTIxng2zKFSVQspdJ+s4l8lPV0Bh+s7qS6nPMJtrTxRTZpW4OPD/5XEUqtZ2hyzhfbgvD19mb
hoTypO/eWaLHOGwwVySiBWJRmkRnf0q9b4po8cVlwFL0dt0zsEtSlt/ZgneQB8yAwNsF6K7Z3q01
ruade8o988C+gy7/X9MoqWXlig9uIQ0HeBSZ47+uQABHQdG0gAUo2G81xziwU/ed1zWDenzlP2Cn
Rzz9pl11jsLwiV7aQuuCqPJxN96BkB0Yji4sami3DYnbzyBP1oRsxMjKrCwKvkZZ/se1ess0dFan
fKjJOD3PcmQTFpAIqg54SSVvztnG/zgTgz0YUga0llO8jJud9bXIvxUD069Jp5xd5bt092aagzb+
7/Uk3BOWW+h7bx2Bf+BIbF39yHezQWJ8qcfbTHyVuw+cC/ae65LdZOhM3MuVUd+sdRPAJIg2IKf2
USlZQbfCw+Dlrs5Mwv8Jzt+ETb47UlylUBOXYkpNUzQTeYIMJuVon4pFV1ILF7GFrk797Cw3plyS
7JJbwBsqxI2tGKsQv2BBZiEKfuYljLJqvweG83MAgecu1aF+D5eEJrR7azwtYtJOxjvVx/VlR1qf
Idb0VGN8Jhbx6GnBb6yQwA/e3a8rFUDK52+tTDKbhFmb0zKRejv3CPkNOq3MdBQhwhNE0ihNbVNV
adcyPHDa125fXHWujUUM0k9EdfW4vhknDgE2oGMO40xsoIrelYuSdyfAzlYMF6nNVO7tYGOeGBVD
WqlByKXkuKJX4tRYKMhxxoe8h4R43ejCs8TrfbsEYnS74334htWeDANBOYtHXKlW3envs4Qqwiy7
5QGHG8yacF/GUkTs3WhCmme0ZtDh8H79/7px/0hCrclWcWfnu338Yc0FdetvsAh+J/EYbgALc2ms
y2G3HbWjIl6y147dvAbe7BKydYngBjPLM1F3IPbdZYvyVtNpc/ai2OcfORozlRJwb04ytqLjEvhA
J29XW2s/9E109JPEktOUK38cJ5/2eZprRSStRy72ScwbPJBJwsL7o5zTD6xwRHCriXQe38GwCHUG
gobyrg7JOb00lLLF82xpjF6cY5OoH1J3De80ZDEjYtDl04G0FzVMsHtcKTfg/AEJ/eWQ+qiOQRt3
NqZCUUVdnQqyH6nVuaQWAHiav2GuOIKX+opUhQY+aB2CBAAOkGH7NkveJ9WNzhwbLxp86LB2tEHS
KP38GmtBAKMRrrEPvT5KZ73o/MadEDTBpbKRFeQ55ofd2qK2HvJKxfUxJvkv9JnWQvF5YCvNf+yu
OhlQ6sh14INoavkMzcHZadz0SU3BIryHktowq2bEuV4IB+ltDsd4DzVUzuRpMTBg2d5CCnRynSgB
OCe7slgJy1T1IqiUQoL6CfLN5h0pvh0ioxXpArCbgDLWXqIIu2gJwYTgU9C+k8+479EEjZM3/YSb
OFe29PdHqTfQiDS8MOwLPr9iHBNwBxGGkTTorGJqS0Qa+lUFxQS+pORsv5cjj8JFMX4KsC7jmjls
kWl+JEAtkkaxWUxD6GrBn3s7Ke5LDiCVYg4lCCiX2jXYGiH01DSpK4KSeUPXQuptHBh315xPUHBg
sktAOeBw/5xVO2uOhIh2yFDmPFCYiX5Ba75w7mhV3Lh7KqHERbzhDIQR1mgU79WkDkFY2zp3VlS0
kRuUiNzi34ppTTy76vPvyj/7lHhVCVA3HVL0U86Rs7a9ApX0JEY187noUAO8WdHxIreE980Y2lSK
DcBJfPEyeSrz5O8HMCt2ia9zN3cWkVd/mBdGuTl0t0/s4T5nKc1hevzb65H9QrYZ9ylYbVbFL/HW
12ttnjky21UFfsBvAPNzqK8kqaFNmwtdlktQxUXWryuj1NQI/prOuXXyg34g+YqAocokgFvcgzsJ
EcqiiQw1Lk7t/QaSozRaqZeVIvAngmpd7z5XlbIRTGXDYR5xQDOk/fJQhaKjdpNoHTygtzNL/vdB
UKoX2vp/973+KdcvNJkx2bbOgJYAM1XoxG/KLJ0Bm/N3gb4XpVvJi3LusTVUGzSfGAj+IevD24JB
2xFPK3sNjsYYBPuht/ntDwTfHeChHANbPxtPEmDCbFwanXOWz7SZIl1iNUMZhGda2zwwVeR9rk9i
35OQbwSB+N4JJn93J8bVY6tEbGMV1AvUKNoR2X/JevocuE9R4Sgs/Bfl90hI9VTiUYmrqqh/TA4M
5xWghWWJGTatQj92Xp+tpRn6VFD3JE1110GWFMSiAErEzEbfFY+RbXPG28q2oO9L6EkLh/z/OWfV
WEqhDrn2BP647WDGAabuhSIXM9DvlJ+uWisFzgo2cQTTDvTaZZaayZ9nT9YylaIfwW3KLfuU5U2l
+d/HXNEkT8qveR6WCXrc8tRdF6NnAaMzjeuQpBqlEU8lhma6iKKK/xe/3VnlmNuyynm0W6E6jnVd
5GfEQHsJHGseNNgPCkpMneKTVRilHIJNihu3wl1J44L6lFw4PS7LVkJBPgVi/AMobtOG2gyCobVq
neOc3/96AVNPutVrWId6/raJDDhAJ0YNEqfxUyJcSnqydjohLXogL1zzEFOLc4WhjrvJgmI6GRpu
1PjAhIj/zqKPaLbq2ugGf0iMmieytAILAKYd8cECDy+x9PFjCG8cUDWqFlIPEBuWqLuTBenBPGTS
/7ocZrr6SRRdYI3c4iJjB2hyFhSN5UOHzYHjOSIzFSab9nS5eGfpNXwxXfjsr8CBBAjvxjZz8PmO
p1BnxAhxwokAu4eMhj4gsQfd8bIIeF3IbduefJZQOrp1Y9UvPkrWv1bcvtTs9XcQZ/UXhWhbkfBY
8Eu1tZH4yBQZ33kTH3s0lbFDfzsDWypP5dovORl2FD0Xgn0aZIqCeqZp0DVF1qWfNsPyFuVewX5Q
nNqD3n0I8pU39IzEflOaj9sX599Dg6BmCkExMmpFXjBcpPKKb4jfJtizlMww33oe+ZVzaYbpk2hc
qokbZTdBGsT4C+A7rTIZL40msYrhDGeQCttwTm50JN9cRRL2jKWka7bzETUpemqiZLe6DP1igJkB
TajMqYMmZxub4rMes+lqw8SI1SqeDBClvlU2F/GPlvxzauKt3wJBsVpbiz1pvAFpuH6AZM/Pi/pT
nGBrWslGLm6ISvs+uSzLWGvfBrlLmjWr/SwZxZTIHgaDTEuM2dJbyEnrlc8xUjJAEc813uS/TxRt
CVazGgfmVtg00ik2qPf++GihGIv/YZ7WUxEsE9IF2MCc/GSuinQ1L+csLf07nTZMh55KY0e2uIoT
pxw/kSDoFWa4jKeRwxkJkHiuFmn2chj7x8dr1A4zjT2KtMiInzvUVuVA+o8jsMy6JqyEJFJXX1z/
1yOFHlXLACkO4g6xwmS0soMioSNJfw75Xg/ZU2zaXhDBffIETcIblcUEqPlvGUlaMsXjKhxuwShY
WVXHwwK7AE1g3gu/Ffd13VmmcGjapimM8rOCeWiq9D/w
`protect end_protected
