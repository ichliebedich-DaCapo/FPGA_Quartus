-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lXlgxby4jACFDN8g/8tgTaSEHrKb8cNSjG/xNIdykJkPRzNsM5TfwCZ1D5IENzPD2aLsSZQ4iwdd
YEopQ+3xRlNCPWbAiw3RImfHu5UjF96cCAxkW9HUOggO6Qt3RofNrK3HhdN0NpuC3I2fylYIgP0G
r5Zh0jLfN4s92Jc4StU6g3nkhqnGCDxteRfBxiftbc6I86lPijEhuLe4bvCkE9GJv/qQUJ52ao/c
43MTqAkbw4XIekQNuOfD7jwd0IsjDSRUGL/GX7aX6DmojIDGGMYrbI9eu8sh/hIWI7KpgrYjaqyA
68L34/F3NDaTv0hd+8qIyGZwHiglvIck2/dZZA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20736)
`protect data_block
UdHBUdaUrQg458UIrjMaq6d8X7gNBmir7fcKMmjQv1Ql1KPTeRQJ854MpN/JrxnyNLEczjlrnF6b
/hkvdQtUnUqwU9axKEerhrn9pQ78jvLIcSPFQlUy9gBGb3d4C6+C0dNrYmgvLD/mSVEb72ENvXdr
4Ap6p4TiLwtaGVQUd/XRefqsIkC5FojPKpg4NCq/71gNyh0Dk5AMmFIVQup6kfgT65T/2NVju0FJ
sXl+DyJgIEB/y0Ok3kxnu0xtmAQw0iDciLy3BXRyt4gvyio8+pXQ1iQvXFL/3V7n2X1Xo5otFPDe
bpI100Nlwc9sCbu/GGu0WXM2RswNCETT7DUkYGla2Gz9CC6EEAErEUr8So9nmZmvd3s3hHaO7mP3
fEKrAMVU0ZfpOxFGlCUhjZlw3ZNIEPZzOL9SOkKMvsup1EvnJHa8jzldr/tpEvYTH8btdowNsNkd
xc1xmIOl2I90XwuUJf27JST+kazo/w7ZzfhJvbzpk11tIA/lIIGVMh1cQCIIYw5PInBe9zOUgXfY
Wnr4Z+3kUIhMOJfjB/dy6VNOdezktPHfEXlHibJThReStlggjez1s9xlnJ2qYZbsiP3SqPNKp6GQ
ogDCU8Mpivg81focUtEh+c+ETehe3OxBLUHCwITQ8jNaQhjQl+/J1qtaRuMVxpA7SpD2RWl9jBuQ
VMobrK3ppm8p5ZJqOx8UC70Bv15eHWeBAR5+GGFvOI8ouiaHzlqGwJMJlLdZlG06p/S6iTOjPWoD
euUnyO3aHE95Kg1/PE5ULjw5zx4TScdi2pDlMHmwGhtwJVd1cuLMC0sVRRs/RsskY5knEiG0abX1
g3m6RGwA+TwaNFUmbm4AAg+hA+iv0YPIZPfKyUHS83et8J5i8Ovul6ktyu0e55EynPp3xZx6I1xb
gnfEv+zKIDpFp6fSZPXSulXfUy+55hmliyTCtn+YDQDUaxqVMvXiRs67o+wQyW8ogFGD0/beh4J5
FbIdLwqIqAKStEcW1KzKUnMhekuv3E/BMLnhgkZ4sgasbwzRSnhXH/62JaXlB6/mYnV8SZHrU3GP
PE0TC+UFushz/2ZSgZ99Pt4TI+RgJZxkLzdwCJawXxExSSL8SK5RSAi5GiJYdzUeztUnWLVPzr5T
0PukaSvQUrxp+WrEEQzedHtGvmCw3hhJNQKmvwrRs5AK+beeIGw7jKxpFh/gxrQj/ZgjKxoeU5zs
JibR4R03LJU3Kb74UqIw7DwmRv2yXkd7yj5YmVxprgEFYRi13wtKHD0iRRtSKW2X0RrrfcEMJvyi
LjWDY9Irw1FCNOytF3TeHVXlczt5nteE5+cdSDKFpgr4+r4s3pBDYQlwzTl/5Bdo1z6Hj2dSEfgK
kEYHg4l9woa7gm2uyIw+p/Bkdetss1L2R6zYpFF0AYLymY6D/UEY3e4rDyLdNVq/jC1Gd5C99uku
SUA+md2xgPasLl0Il/60SH7IdNvnwAGxjzkLeLfRN6NLakZmqP4GipTeflxi6UI1nHixr9rjPU6N
YQgkYj7bVuVUKus/PpcIUYCEJ8Azg811lwMaS89+3Od9c1qoA/92x3NaAs6ozuXG8LbBl1x6CHZ+
gPuNQpwIGSktsJNsZVE9awuUIfLRZYbia/6vM/W8UQnMbMEN4PyBRDthSnuJQHyaB5P+Az1XCXIh
I1DzAX6SRvGvyeD/GNBtTzGr0d+tzswOpVMtV+69VTZfha4+VBMePOCMs7Tumu1WqZlsbepph35+
L2mdATOYkzORRitHq+0VjjG/l8YjfPrldxF+QZwNRB91Iq5JZipfo3CuCxepvu8MmGHgbdqKd+WY
RjIpwLE96tcAmQe0GowwZl2nxDd0iIgq11uwMwe6YB4Zmu5PiPaTCWWvUxiLTXmFY+7c7Gvyym1o
afSF152j9X3z4uiIIBbqR3QufOsrysdM+GXuFJHqAQ38hYYiaEdAx10RE45Gi9+eZPHa8BDkAZMy
+7i1MWkFR0MHr2Pp/Bo0VVfKHBMiYRpQGEkWqX33nqdNBPfFSBTy46U1mL9YOEcYURI3pyvGBs6n
lKA3jRLQ73klX2WAijwbXz18vbM9k8m2WvHNN2IIkZ9t9RMYv4yKME6/Gi32Sl3PqXRnfeFQyOcv
bUQC7gj+YjpbWCqXmTCjqLHWJGNI2kD4VzVKIHmVNPHxM5OgNIpV2soaoNNd6d8lzq8el5pth3BZ
Ql0CBTQMdJuyWKjkR6i/IWEaBgCymZGngfp9YT1bQO+uOuRlQqwnzyykVcksbBWojqjHYcITcW4k
cTJPgfD0F+35Msxta9DZ5PpxgvsHTxgPbFY5N0nFDr7q8BxvnbONFtqq8TbGt5JKPQX8GTtHwcur
EqBV7TVi6EBahRbwh4A60RnLCOQ29YJzOeNxPEbPysoaMqzIQdYixKRB4IPiWQ3tW6TbQMw9zFR2
nlLu989zZLnAYVbeHWAG9J7s3tLIygk14HduJeZpGLN86+X0YG7PzNMDlgXlwvNpMVufO51RP7tL
vu0lXhMeTJcstd+XpxxQlnj1d2UHYSTT6Tfi+Tk6wHAGTvcnvnOKpnJ5SaZz08jLlfstmsJSUJZh
LrPbiKR51SvrJ1Jc+7Ng+m9hUxi535RVZCIy9tquu4LK4XwP7CkOULoLDOaw2U2nR1yfR+/qDS/H
TN472qFFU6pc0zUyH9INHUb49Y3sYafuJjdrtBkOv1OPPrU/M+G8h2gFW1x8NBy7k9u6zCUlqLjL
gxD6xdAbY+/8jF+mWNmPHo7jAQS878k/j77g7ipIH2t0XLU+/7T4Rxj153jfs/2cXkYRG5EgGe17
kaXCpwDhE9/zJERZfGUypDFYPTXPai6hrlWpr03trw8GdxuH1u1fWv2qGm8f+wPPOaCQSoV7akNS
c/qPcT1DRchvNrQQDAoDvSFPu2j24yfLhR1Hydy4OsGMkCDh0VzQUMC3j8U48tPVieQusgBFw7kc
+zTvym5H27/VezX7HpgiGsZqLVqTBg5403yT47Gu4xCLoQJd5Z03M2jWpQ5SuVAZO8KWhTalU507
VViwYnMRkEvHS8C7YN0M7fO2DKEq8M1NxsEtmVvHZBXMJeIgzrGohnHDwD5S4tnyl4fbHNVgUNXR
iL7qgMufKEaH7x/JabBmNXoJubv+COhGJCNk3Fci/uaC0IBXMUTxdFfz0HpYNnnPB4FjoWQBvDDE
/ur/ZCaRtaA3rZJu71bHUTBJrHt+TAiUYjiNLOl04cCd6MrekKBjYWorArGYHQmDxem+AQpR1zzP
bC7NYgjav3nqs5zFvfzgUKAxiSzfIKBdsUcUWwNtzklFu3RCo0Ng9RGhRcV18txO4sgvEwxAgoPY
+Qq/BLhndQg9c7ob+kkt+8Xv7umhfChCnkMBLgB6MFrmhf0aCTf5TcMvlxA5QaHzQBDJCRl27F/d
RjCsfXnMHnNeognrXDuz3hPfvS2b5bpvdyn4fkkKp3+kzyKyfwmmhhbnhRdWNY5sxh4Pev60GDAk
IxUgizx+92rrwWCJ2W/nytF6mHVuuuviYhikf+9ZnCXrAhk4Oor119y8UpaYSc5bdi++h+1jiU4n
sBwSE2JRDm1lHveCT7od2ksDd1IBD4J4CnYy0Ta03OxI6afKZ5lPr0oo0G7F8G0a6a+q36EP/9zj
PFo3w9yhoi9A8BCpkA29O2hRWq+H74od4a2rXF22CcLZooZAvhYXecMGf1Kd7CWbb8EBWzNuK2yl
wXcTNJAZeMKKKhG2T118cS7pbv6HwPQc8genTfN+SpteW6SS33R3RVKhm4c+Y8YmBbl0KYnbNqxi
GLr4AaBCI8kY9YIFsJI2s5MXSCKJOU1TDFeRg/j+nrtPvy7Rq1/CSBRTM8EYlGpZg79PzXlWRKd0
BFAmr8fuSruJbaDOKe0clFdBzr8mXN8AKWBvoCq4BLh9W2flNmWHDZrrJj3GdaYIJP8n2uZNv1fz
ggRLdheZhwDKdI6bhgX3qqsEmPRnYIlm62vH2PjsmhhPC/V0PqFAU9CWyMnsOMVNo0jk5oraGugR
R16nIVnz0ksbYg3hGb5hJWh2AF8iSi9yx2A2ZWYeuz5AhHHk9UsiAzzYRttGf64BYeerH4ZK9tVN
mf47Kf96hJ//Athn3yrNXGRB7FVDwxQSfnRagFtyJ7AbTtpAcSdLIfdcPMYpIuQTmNq1Ldch1Fyi
z3vip8Ot+ZbT3i1iY6hSGm7R+I1L175Rao8p7fXC6xt1PyYkpWSIsSa059sVbIDKhkB+pCGc2egw
AVuoWDi7J6M9Fq/M5F5d1MINWV8QOnuhY93u8RE+2kfDg8dXJa8RMdaIOa8JQ8ppzjF6AWROB9c2
GGwYm1Ssy8HWKW2CcsGu0ynAz6fsvMMSEgaA2IL554qW6IRiqimifOhq5FoSA0WQ8kwDOldYxhcR
r/B+7r0+hSC8+I7w76CG1aHJbWSGTuFIcHUMGlSQhNHXBBuAdRmsBnszG3vWJVVNuVVH24IeZ+22
CVm7x+WfGugtm0J3penIriwNZ+esdKqd3vWmjmurJKqTzEmOIqf4SiodSMaCGHscOv1jfUJEGUiv
brxqq9cy2Gfe9hNyOTB0nY0+hW5zKn87XS0IeTbm8VCkySWeYJFnImN05RDtpPdazC34G4KWVlkH
BrVSc1nNNOGOASj+XbIWA2mcdzP1r3OsRStbQPmn7SiXLBC7VoVDIKM318qhgRk6mVoGh7qYUTSD
mYOyOs0XC5n4Nk25DKppgzwAocK6IMPIliUFUWmGtx8DBiqUx5GZed0EO/4+1a6PrUxzjuy3viLy
t/Ift1fOxS+R7IKNrvuJexTySCmyhOYqD4MgDEBnRFqVWgI8lVQXT5gMK/dNRv2zTPSi8UuvtQGX
dOf/lzO8H9T8aEA2L8ndzQ+oT4d3cqhDzVAJxa16X3VDdqPOE2RBnUXJNRB7Y7PuudzWhP3GCXOy
GA1JrAn3QgUpaXGVFk3Nm3C5Arnus5/3PTJS/e4WtGB4d9VdoWSVvjv+3Xy22VK1nsH0wnutI7x7
FgvkUFQYykDS7cPjAs7AuDlVVZxAP1HIcNtUrIlfn+lTPSgNnHBxIeK+DSNqcQaNtb3IkJak5p06
iUBtqMRdBL1ECBdnrU8lblh2MA0kVUc2URfOoENNuES5L3HV9PSBIu1REMIozUm16A6Ukh8wDJBB
ONTQmJMyRW5Z8zrSIS8OholsMWNEhmNBXpNzc6aoB1SM/FJSW6ofFznybk1dMA8DMRGWJV4Y2n9H
anBeLDuFw0Hegf13nHpLzdiNuZaZKcvh/WGZN/xP17wNgEurrO9WcKniGgXqxyIgp1zZsGUlovSE
M4pRjPlcxk1SuIClKLSna6ANq1Ix1Oe80pASpNnYZFVxiNteUTOJn/4E8kCRAE82Ni4mScQd7m9X
vTtPi0lKGdfTd4S9LBc/QabhYNI/UpOkjNIsZipRi8/jXtvHd7rOmyWvL/6qxMZfK5GpoIKmRfYK
80l4ApLmbuMpQofrkIdnGxLUq1c9txG6/ZM1C6ysya06TL3Nq3dehezvT5ZsajkBxnelE+lW/Df8
cgyI29FtMFH+nMvX65VN1xod0VcEv+2/JpBiNxOXEvh5r8lp53sbTxDbNaQf8E2cLVuDutx+M55Q
qGIGyyVd6VWFf4rNGzQGS7Yq7byKF3H5sCGilo3/LxIVql4Tq3LnQIfH8bbZsdtJ9Jb0znZqHKbm
IGDAsWCQzvOsZ3+Qan9zlapCvUXPsR/rvN3WMJ0pcDMzqGOVTqD+uS34dMvkEcJVOo5YviiFUXpp
u9nfxOkUqNiQXPN/0H7UPi/JPr1RjkUcUdo0MHU93YMm144oc7on53I/PxIgHRb7RrI5mBZvVQUX
Z89JSAMYJT16UiauTlvizJo+3jInV/04XFUDVwvLGo2qGGYEdDPrvmweBnp0XWi6I1+wgO2eYJEV
9cl6jsTxDFFh22mA1qgifEsS2NnWsvkbTg3YKKLK9pT/KTyvezeF7D3fjnexR8or4Ytfhbjd7WQN
BzShZG1ADrDSIn+8XAlt/BGuz3YR2Qy1+MMlSjJKAYpHAkeFAsBin2v7XBvmhm91rrAUfPyV3XQJ
A/d9oEjInn71n+kNlWd8y0MiVpGdkqdnxw7wjSSEwfh1GNlcTqTo8eR7G6c1ohtiB6txfSGjPwtC
iNPK2TpiMPCX6TqaJpS2eCArNscpya7k4+6Dzu8HCY4/75hTNdfy4LMZFPEmCuIaAdHm8cakITWz
5VWbULqfYVL55Ixb2J2svBBIrCgZnrGJ7xD3M/4BmlF0FxbpK2pveQduPLUwRhKtte25YcYxm7ft
nexw4lp+RkjgU8gBddDbUsk3tpX1/exmAqywrV7kl8rmiOtvn6cZw7nRwDb/VPzSCJk19rta2uY9
XrTRUYq+C2b7bPLjHM00C3RMyJMi/kxtHt7h9QDNERNN4uby+41O40DcVf34RpvhFwTx7BDZuIVS
/LcHo0hGWTQV5ltUhcJax5s0uYIfVkCUfInXlxNKkc6Cn5DXy2L8TR4kRe/9T2uTvDilkZYjHOQX
gyYamcaIEu9FCCEQbzOHk0oi4TUFtdJeYz0AuQCLwxUk1PMZJzWff/sQQridSvTbIe2EAFdDdC4l
82kpzwlwZsqLoEbstxzwjoL5S1HEZ51DNGw1nHH19g9jYWFYtpliwSzBh16yWfVWdsx79O/TjQ+L
XW+P3zS3b8eUh4wsSGrounUdE8oXswD2eKiMxtp3aUfejG3kk6g24wxXhxovTlzSF8piK/7flS4d
dh8WGHZtKabFlZ0JLby0pLSE70d0lfJQLZjCYBH/owgnv2iWqEcCpMmn5mOV7+1vTGBhGgSIDbfk
OcyrVe3O32x1R167YXBf6syJvFon7xa800HikVknp1xPtqkGR3xZHtzKwKdlRDESF9cQkTTW3vdC
W+aTHVIWbcGX/4eFk3QA6ZRepR34Tx84dY1v/PMj7fDgN2j5VJgMr/kwwUAOykZRIcwn2bzPA18z
V+vZRw3DpbyW0yOv8ciJ3IhtzDBKDLJrhoWsMe+DDJ4m12luypoPFAa8kFn1nBL8l33N05UsXZsZ
WGvzEQe3hGXze6oEXIBG0gXUoYq/36bBSIOZDUy1LNVqbGJ9yPJkZRZY8ubQTkzYvINSG9SDFY6t
ftnb97+fNANsFAtDxhB3psLYqMk8nemTmS90MrELk3gqHz3iBo+9nD+h6QUG/uUBHZECTpJk8i/0
bFcKVXDW6Jzn/avrZ8f0KN65BxSgwPf4bKYDQpLgmEjSJ91xHDbg7ygoEocUTz+HHhygT5G38wZK
/DeQwlWhF+b/efDj+8WO922807Mvxn88oIjLLmddqWfjvVh9wY+y6Q16FJtv2G14xbdLKcXoFa/e
ohEdYGl3ql0lqnGHdQSIgkxjn3iyNFa1S/5/sP6UYVh30m4lFSOwI8txYIwPlZZtL5r7BSYQs1ws
zNlda0Goys6liqCU/Mm/bw+6vFGLZ803xwkJHo4NjdJGNmYLQrFxiSZHV6Dcxx6aSYLF9//mrqlc
TIlkOLIPINiH9WAjalwMyI++N5I1Cwk7aRaVR1JWDXniC+KZqyGARf62LRfPNknMdFVOy7zBGQmx
CL9/ZaduukZwEAuzfnRWaNV7Tqhd5fUievW+nzvkba69QovsbPBs3LjzWKmjMy4TULMqzeVSfeyt
/A3lNQNxpK3KyxLQKofhilcHadHXSL7df6IrXzh/oktmOZKYqYQC0BWZqF9NESw5/4hA+LmxCkas
z8tF8uTkpn70dXNOsLjGkCNGz4+BTuRxkXJ2YIA9l0aOTU0Rvl5+XhMYu0jGTVe6fis1heQ1NIFy
m48r1dIEg8QUKAj9dR0ghSiYmYxFm7MLZSHpxY/AmkxD7Rc+lEPpRvjyX7ovxlozM638PrcEu5m5
7Ds2ZdbjlKwHNCToDwkF4JTKXnhipkQKSvVvW3MDAaaCVdcX4nlamlzDGulURTAFbzPK7wnnjmvo
qu4IldAHOJ4vAAWx2cKyHzuKxW6Iq1YMJXqI96t581Evdh0NmDEPKODwkCSFdcQYtJ2iPoAojqVw
KWI24RcKsDUlmrUFOdQLR7oP3JbwKzcrqPGdF24QIngVdeURwZVaDqi4UW5LPbz/5ah5WUgi9jtk
03G/45CCkm/WnMUv1DmRsggzRvtYHxIb+LW5yja9rPzsswrsSXLMs6xn5Z0CE/xz/VidcD/vk0vf
5yZdppAo9d7qoBtkPKzKmHzmgV0Ndnx5CDrLKVCYhn2yCxX7mA+BjRVR8brvtEFC8wZAPUwgqrCH
yQWw+ZMI4X3eRlVz49Rc7krMks6EZsXhpmAU1mnRz4P8ByTQZ7aL/clcPj83/Q1xTzr4HE8SF1xM
M2XkZqW5kaN5+0Kxq1a/8JrP5fEL7LaoCWpDAhbmE2NU7RpiXuDRtLHTyGd70kr9EiJhdi0yL4ll
/Kavw2pbBGzhbmbTC70Fe7Cav2F9Z+UQ8R5OiTWEuA1Guq7745dZ9zBUWew7Ragf0z6iQUe+jbz4
ArWZrFHqRnBAPsjkqO5uLbNhfWWqKWPYL3z398BI0ILOQp9AdLiFmeGkHEex9E12z5YsKjv6QqW4
n5mG/OgrVFFzExQ4BWyKr1Wt4iOmAt156vgyGrosXsxD3dc8uplqWeyefOakbM/XyqJD10FXhsH0
hq2utgClsgLpYuYjL+Zlk09tNrHqnOUhzlCLqTSkRhYhkH/A9hSmSEVo7eJI51SEAQfJKMaP86jX
7UW8XNPG5x+2BGS5c7XBdPKSkl+egzFje/7nADjCW2lYOCgYytdclaOalmPksUOJN7VlkbgFq4zT
McnDJnVFvI6aYgomf3r1fGkUPK+ktgaw/NR+nPWc3GQ5Lyi6v8ZRaJ+tbaMasOvE6v+vdyV+KcH+
Wue1Q+1rUnUsY571IrrJ4llfCXuDiwJulfY6YHDRuiQz40izbdY1wdupIIUX8h2p70sV98OePj4M
8Tcp+i1axJy3gFGvusHH3081AsDW5BQdjB2+1tRuAF0yuPTzHwIfzePPsGBst21x+a/8r08bW6nr
uc22tUUo3w1vQL0BCVKqGq96Lf+toNobqLt4PKhlh+3wohHAjZQD/G/hWjP1dTF98fr3Gvglp1yh
HykQEie7FlhnCnLaSpMH4tRGoP4D+/tmeSyG6FYcarSqz2XG0OmclL4OsgdCGNGXTE4GTrEblVhI
rqPSWN4JjPmrT14zzuOdxlUeDwH36GtmcSL9OcOdeQ3azxQAhTXjN7iZmZ0+iGwL4V+SXZXxCq91
FfF54k/FKVigxn8dAWeOpxVJbkPAj+s7PurSfXGOHygstAM6Qdih4rWkA4pm4ygL8DrVLuCutNo/
JlOD6cZ9refKUqKWy1PuiKLv54GUb4hbwOqo4pMtEsMYi7lFuVw7vh90w1h8qyVEZWlU2htKV8F0
AnGmuT2zISOlDA7JH0HQcmdzkGXirIbNAMQi+LYl/oFPzQPN2SKV8PIn68hLRlQ19zMRa8PXaQXo
trgbfHhMLhiw4nzTUcIwN3840bwbgxb4C1W8cbK0U9L/sVXekf1oazKFx2x44NVk1TWQLfEgSw2f
jXqd8CrK0r3iSeE8ZPmeOXL0RBEbPOqDwSUxR/Y5w+qOx1zQSWXCDSUY+uDF698k3hStTTnHXahd
pIw3Cvw0DHFzY7Ww7gZc9uoEaRQ8EuyxJ1Aba46OUzlx/guHiVzplts0GrpOVPKqf8jmqZu5xJ5K
B5OhUT4B9OuWJehicgiodbAlYoLJu70R/b6FlCf3DOhoY1LgJNqRMp+ESvopracoV1TScK0aBQYW
0h7DOg8skOK55G8sCLMvVAG8lyhOBSW3asUvL/dqmMuQFk8SAwVLV0LbnFie6e7lo4cUrpozJOEu
FNqXVzwlM83knYmiz412nkUpmAO2LmVpXdzfIUBUIZR0+QvAnHsG5GWofbgxNG+6utUsG07E51pH
aQ8x4ZRnmkbwfF4LHu9uFHutcYfz9ZNUlb1q8VXSAwxLfPlv21pzFQqTeafaebaRz6kqnLlhcco+
Q13Hkxn3yU5d6NDdTd2aoe9IE1SdNp1GG/Aw3tGeJMCEBbqFDAVv0DJKdphxKUzBCrhs+6/E+GFP
YvvhzHT142jjHmm6IvBHTyLelUUJxldLhQyNufaLhEiBwV3J0p+NsSfLTpV48gW3VL+5nAynVz+c
cxT7Vv72vdrS9uRIbJqSDPO7utrHosmTjwQ/NhNtq3tQkY5f14hq1/LzGcwEwkIY+4DtYCoEs1Gg
jwyzhT7OlHXhcQBwcnTp+qGn3oYos1Yr/bXORyfVLFU3E6munrCC5mS5IHNZNkdYGWAuyUFzD5ci
0JrgP+4125E9/ULdh9x+BLSlFZLNTmpALdMz276d8vhOUez2GrFDucYXxFEOPdBkOsspZu0nY+fv
aSrerhAxBZ5O0107klByVp4CvuolRAlqDTwxhj4OW5nQx5zvQSNHolXr8DVSNlhENjc5mle/Kto2
EdQRNpZ9MigDf5xgrTvzY65tFC7HPYYNrIZ5MYJA1kA2WOLrxBmjEUg/WTqCWe9R3C5TwxAdotok
UFarTheqjoEj1UD+s2Q+/yaYKmd630HugU8ApUF72BBn3lYQ+CqAWQo0Vp7BxHuj/NCXCvgSpVqc
hYEc1x5eQncuCsyNn+Vbj2PTZ1x9IUChoicpZ7IVdw5GlxLtdHjxRGzCkmfCjDPpzS9mEhux37El
flTefiX85rR/EgoJGJxaAIvCupAgZW/vVdxnR9CmRJBenTTJ2pZY9kxlmnBsQRtHV0a7mnngnBxq
MX4Pnu7IsU+Ikl1By12C8ETL4jGJcSg9D1zy6ZwuxPlkBuBU1zJ2KOUGCnrii0D/KhyM/7RjOh1d
VHZ88dxbiY1myvFCo1MtcXMQlcWKSfJdyeCBDlXqta5z6x2UW8BKK5CglvNjEIqrLm+Rd672qWe2
7l4+9yqsoy8suVBUErlgz+tonVNLcnRvyIJ7t5hul4lfsaLzUUV2xAGYu2ALX1P5v+D2r+ZALrkq
9coEB+KjGmbcQPSWbxGMFi6ob6RG7s+R528nhyeVzQZWRggHzmeRV+yYQsduJfmFnD01026u5FdO
6ii2UPXkIFTYPDuT/YHNEfr5FlATpCmcW7zqdFz47BKWIEV5txrjFUO9tG6369oP9JQqbo95Gonn
F1pwGIpEvB9muyE/dvmJOezRNpJnACJutQIpBHl4MLpustYvhzB+keeibhmDP9UNyjzL3i9f07MZ
BRmBKkqQRv+jryx1vcoTOq3s5RQvyKzpHJMpPSpD7OPv8zmMwP/uNYBt4ajA/OYmA/aQtQlQa7iB
FDbZJUDPrjVIZPrj2TM0WPDBD0EjgkL1WqB7K79cHJU2+0BBlnrTkROeorjPE79vpv/rixt/pJby
hMoStdmRHPniyzc/S+eZBXOvfO6czNmLYOkpJgKARylJOCiIsF11O/moHPWqodkNgo3G6g+199Uz
eh/gC+T0zdIuA0UNOMenTlSwIbt7gPHAUdsgRMjhSqxhIdZn/3wvez2O3urlxUOrE/j4jHisPF3w
WXgEOTk6NtzTB2T1oMsOYZi5YHWYrgEODF5oQaqMkVAmYFG/KT3At31ZPJDtr1ML65sgFJpG5uGF
iNhxGAXdTucqIYyN7oow+vnQAnNeQfTL98o25t1fKpcMUiqGsOZWmKYeVRFBnp4M2t+QauJ/Z63O
9Zaov1y+JsvCyePgdLLXUdSpIy8Y7sUOwr+cty462fARRnc2MyuxIguWPbATl4MHas/dXJLDR2Aj
A5U2xU2SAur9i27m8Hga54KwApnm5cBNa9KXHGzICeLopnujLFHVLKpYIwqSJmrn/CNtUKenpt2S
bRAaQK3aEV3v0cr0lHP8Rk9+x6oy59rVdC97MBesyLEm4ReKgAzkTFL39G6+kP9BQxqruWKypiEF
l6hOYmKlZxkY9FLtlsdY7XO7pbG1SDuPYyhDpjj39R+lxFPOgg9EKidSZlSVYbxfY9MlNd/CcZGE
nT9ThhUGw8/57rFrBXw4jBanMEdhtpO5p9a4m3iut0J0gDz2cIUQ14exNA+zLKqulh2N2iUaA3nm
+t9DEVMdgrxnvyrcY4e6WWw+IeFV7Li886UBSv5b5bCj/fMjGZnw7yRbvwT0DVEU2ok3UDyb3+7n
WXJArHkKMHAEze3sPuQ5qEwIFBt7U7UWY4UTlOzIbTULmbkI5loLHjSroZ6U/HxHduppzBYe1+M+
yq+tl/U3zERMFbgTFBJ1+I2W/TMuTVqjTdBn89tN5hCYafQ+J+AoVjVQFq9P7S0dkBGjVgyTKSOp
eG9Q30E8XMaoF6IrRit9znon+dwPSND9kiePz+YN6whOjh8zNUImgC2vb3EYOkDrhu0AM1M8UOnb
O5ps5lFCYLIdZ/Vc0hvBPySc40rHf0DNennIFkosQUEmTZmlRolaT+GqtHLzlhbioVjMh7DG8D1Q
2+EniP3X7kG/RsYfCEdYUg0Vh+krUAwc38UTtaaW7l9ycWkvKJOtx7Mqq0Vux05+WhSusipcCGTr
y5/vEvNxJdU9IJscmrE1slR8epaoyWR5SL9lQsNRogyXMY2Hi+ZUfC+P08KYK2DLhJ9S3j0ogPxt
U6yXegyQfAvBiFmDPRgXKxcpC8PyjIoEYh/sDhGq1Qt9TNM3CtpOjIYw2wd2Xwcyrz/GV8/Xhkvs
HkL7/29Ryetdqf0AMxyIsburEd32xrTXQVAa/n3CZZCs9C5idx3kFIwQnLPCDy3pExJ6+mVgA5TM
ixeBaq0U3+2vBRpsMVIzvVBbwnZucyr1XfYyFjSHTAe153f8At2+/Qlnf+Rh/jmj95PwyQD6KfOX
mUTbt37suv5xeiHiCBZigOfDqJxjhdsYwopfFWboLlLxAWKWOoYM1mY73DEkxmqktdED0dT2Y2Da
Xta4bXOiynbiAOuyRKo4VR3YfsuwBnoiQV0CLmw8KFeEE2erpwSUwfE+8YbONOnSLS/OS5uijhlD
FDVsA5D0cmvrddnbTWhDo/hYVQ127w8+7SMFnUGf/UoHDM8C/tzC4CKytFcexov0lnbyVRVoLzIV
7vcvoq7XE6v+avJQgl0ONz7R4h1pcTPpMY/Hdb50aXBZw1rI/eYCEtpB0x4862oTX2ydtATrdLC/
krHLgBgp8T3pHxdMYC5vP2WCk+7J5HeKbXOOSQEjEfxbCPc6NZnKMLkwnSgMMWn3ESJvbmf8Qcr2
cFfyb9y0kv/0a7j8ly0iDsiP4vnsOJtxVLmFyMaEkSRY3dnUk1hq1GB/Mwfc385HrcTBI13fe9rv
qU1txUvnYHUaEGpdtuQbzZ33nl2tyVdtjv+CreYAIBuIYM8usVQ6XxPeRoAFl8k7vowXz4afXq4d
nq+OecAcpUX+kN6lX/QSVm0oaO3X4owqZVIFDhyFUZaNJJAhLvzHR6BhNrT2415OjJAhfe1+oRem
E3gm/FmCoNn4ojRAnxosiNpnRj+RGMVO/TEwC9m6i8q8sfP6KbtYDFudmmI0wqkyeZusv32HN7M5
fFDm6n7kU8CEbYK+D4BkLI6I8qhDvG3fpj4flCOBv5Yt5//MrZdFn7P2OuqSZHI49aBsZOZF4hMQ
Whr0Ql1q9uAtwYBxTGE3fUCkXzPaPhX0hc5g0Qo6cp1+8xNQAX+ra9lvnP99YO/gPrwzL7W/X/KU
3HnCXG1GdjblpNp9opmJoaDxxRST4+7/4WdGPNuBRRb9G4TUByW6oO5l9Ciuc3nf9h4cQgqAV9qe
gatZi1+9sosZONT27o4ZTyidfQoxwbqMg7KdM+O/hkXyp58IfTZA7SbZRlARusJa7x1UrzrjapWl
oaiZ2tA1Ku05KWabH4LqdVs1+ei8F2+C6A0UqCTTLerfuKDciQC1dGQCQFNQO2nxH8UPhZNi0vDn
IEuO2glTPthDXmEsesnOYrC8K2jFLmR5BAmOBZJN9iyfFn9M9kJRRg1iBTs4ThYTuySEaWcZUqZb
CF6CSwstwTI13HKbWe+IrOAP3ELhfe0pV54k6PteucawH+nYEFSvwImTd7bYBufV2tQEsLbkpD4q
C1u4QjqXojqKwTRJ7w2hKPCK4bxCZss7wr+PnHTQfdjI5uoUDeoV9WNWvxYsbNzMDchZcoNOqJTq
7qG9CDbk3WVUyzks7a0ElojTvNzyMGDXSj+fMh9pzPxrIGBAIJMyY6o0XYkAB1dR0r18ILRBKyvx
3a40LUI+Vi3Ai/7HfZYQfLU0qFgLjk0aSYXi+8i5B7lhSeMvwUuyr1CmlWMKb2QJobRgHJIfjH2z
BAchO6TfQ0zXswRdlVnvZEKyeFu7bHpvg1sAtukNEMz6IvUb9v8ZCXrm32y74KAMaVpJ6VMYiZYL
c65y7fKRYvExZpHYTtt9+yxu4p4ncpuT15KJ5DY1aDxatoW3JjLD5DypI11tSHz0pqQ9bnMKNL+T
nJr/oUaTjyVexvKOob9q5KmOuGGAgg44buPrd1TcTbdVsTg9g6eHXHRrDS/ow0r9Nncx/jYaGdBb
/xgB0NqS6VSs9XWX8ALpQ13WmGTfxH/Xv89QgvTqC+6bfdTY4anyP4repPKatnLJC/uNjco3ksHG
+u7W6caak1WskwurZ8oVawAzGjFzptdCKHAYXNT5vmEbV98euPlSnj6fw/cxZK/Dh5xbk9vwGGSy
QHya9uShjrP/XtM+x020PTCuSwFP4A0PnWU4v+sF56UW/1+n0WjPB7b8qj+8NmPR56X894h1tOu0
iHB/iglxpHk0MERSz4mM+Ii4tOhjqsuQZElbqgZt1Dzq7kAxMScf76qxmxJ+sgI0QCWc8Jb7AJZm
nyxdviR0CBRfr/Pr07w+k8JTxfI/H3jnz4TMoSh3Y00HgSmaT7vvbAbBxi6usgN1nfTvqh87rEoQ
ov/JfEEWdvHHIqR19T4D7b5G1pRJRn0NMe96qYmvuwQh/yT6nTD2bTH77auoM5MfO6jXJmSADHvX
gcyJQIGO0yOBiJn+y5Ph8C8Pj2XNgYse7kQCYuMNyiWAptV1O688lUkFBMTwbrN3LMRehXc2OoTc
4E2Kc7xFrVgYMwIZdB8NdJhtnSOuxSNqiTLS43Wyrw+qMIBftuPwT7DmbAn5xDi/PNIehkXjrGwX
Em7/Oil7P689YG/LiQIAOCZa1BpNClrec7rOiQtpTDicCotEK/qfrUYnAEND07HVlWClVIW4WjTD
BUSC/dozg1mgoleZOWtM8ohGsIZqCxWLTKb7pIfcQqOJgYHAOnbCFDNOcz0D1b1Z94Sfoo9hB/BO
IraqYRjS1eR1ZwX2LMO0yavfTD78TYgDb+7A9olA6rludd2RZRtnmtfenUWh6w1YT4wnEqYSb4r0
qPKbTnySF1G2rN+apGX7NFC1EgbNIU24J+DGB25N3lEHMaKVZ/ADFXB5N5wh+0ceKs7Rjh6iIXzQ
H6iX9F6Wk5/lFdrW+8davHgGDc8xI8CxlPMbAHl9a6Z4CXuh4lkwOozj7JIjJZH6fSm0iQO9yAHF
2RAvneoggqSVzVIH7PwAv0QQtJteimDC6IzTzwJW6GVc5K+jzN8L2jhbOvjV6215hxImgQX0J2ed
2Pw0Ek8JuO3RdeNsYkM8jZzJbLlGDz/T5p+vTgcMcmHFHPQL9k97G8ro+aP4nr2INS6XNlvGCdft
oY9EZb67gR+53+ScjdY7bTKOyrXkIj9iTYRqHYPpDJQV11A1/+hMwgPdWYrztCdg1ItVsoiX9v8I
UKvmYQYOYM/Kubwl3SyD877sNKG9TIa3k+IPduxBquwvqyJD6fDESjMymONy3oZV0bhE117eKw4c
ja82jP7PYADMYmDUjT5i+yJQF3a/RqKmLiZy0+rq1GlXrFr823junu7cg88vHJdSZ6HH1ZsVYqtg
fawsLp8ClnPsPV25GobAOoS190ercnCKjm/IJaqexKsM8CqugkuiEpB/ocHRgwRfl1xzLN34urZv
9LwwxhZv83rQBNnRaWCtkjI2FDO4U3BSQA3DLj0A6lAeH5E8JHg0Rz86P8a8LS74yG+8vK++sD1D
10sy4JoqAvD0etrUJsnIU4tZpnt18wgiN4l6walMtPyTbJnp5inUJRDUl+mRQGoga87toCjAO4zK
/5IOnvWvNsu2fE+TWiPA/87/PND4qEYYW6/CLhEH9nFka8cEWuG+XIdF6eHNSOaSQE/X7vaN8CCC
q+RYeCOf/OkjeE3ZJ+LKup6GH0clMRdxDHYSpjRd4Zsuh36o0IjZ5PCrDwrvOZ+5b2/n4NScYBrb
eBluAfT/HD+7NNWG1D4zI+ejA/ik8d1lJ6YD14OF6ehlf9u0wXRWiXK+cqYc+0DuHpaGGVOmPmU3
eKXZNXlDphjapAPSIeYSBQhdEnUXcsNX+SK8vUWXdxHiMCxKezNb0Dr5QyGfwN1bjBmY6YWdKSlN
sf69PLAK6yhMVEfadGdMLkRj92mbhdRYOzDOKTODP7rm68EmdYT5qkK5/jzmVud9lKI6W2LD6VcL
VPO8YIJ+ET/QYMkxbljeFAkvrSSuyVmJtuYm7djy5zXQYjq1ColgX2mbY7DDu/Tt+G6UaIcuQocW
CQT/mxcc0KSddr7c4HkOK/mWgJOE1OEcwc2tkMhuKyDlvj2RHUG9Sr14soWvTSierQD2LveBttAi
Fr4MWNfkGb0/KbqJAt81cTCZA7wFjQoLRjCvHNs1WW28lsHDCEkwbFss01etu9iu9H4fEf0vkoO3
cBbalOly6a02iKKzswxUoHx9axkRJGW33Kb9LQSGxO5yavkJl9gviFQsrG4XuDKBxpaQjRemkEit
fIOLAUVXx22p/NU9z9pwRb552PI/qXM/DSoiIuYs/3wW6NUERtSwznCIh9UyorrbNgAlK5NZAHH/
heVMcAAISp3mPW2K4noJZwBD180bW2XkgyfIw52jn28S2iq8qSOGtQJEHaapL+xm+VuRudrT9uPV
izAol0ek3JOqEEr5mxhmCYG/HMQjtJAD8F5TYrFLxswclVClOFIdA2ZG7AW42PmfQccO7mfpzrJa
3ocZ69O561bBU+NZOZYqCO0Pqwp6ou9JhaGNm3ZI3/Gy8vkR08gzyJOoWDhfPTIeUIu8PEzeEhwA
JynPltVgQpY02U9fgCSwwWhpTFuuQTWF5VHMhRRjWVPxZe6XIIBMtezkcfvkp5SKTmr8NcyvhEZN
fkrD6W5BLPAjSo8QaYKD0olHAMnPrDQY/3W3KFe30X63pW7liSjjzubfpMD99Y3RJ7jjJRMsUUoL
tqZplJugjeFF7iFtih1xP7t6qZ31g5szOR2tc652Mn6lMg9TTpsJerXcHcUxUj3qlFBrJL6RlSAW
69LCrU/wnLhBn4tqR0NNtebespgzLku2fLkc/2izrq+riJCzAMGdaBvRzL3oBjOe/kWoHjVzt3sr
bZpoXMq0gRymJ35u8/wZon7dGNPCRgVMvhZkqcg9wbN9nQgDp+RPMTxS3Mcz+macWtiRGt8sBz1l
N5EHd/8KH0GfQ2kV6ZDjHcxGyJwUn9jX+aG+VSOlohI4tw1O6r01wqF47PMD3KMne37TClMgK8nh
hrHcX+ygtTcbQoRefBS1x4KFmf0GylHdFS75hZHkW4eftAVruJ0MJ0Obcj9cNS7ewGLCLb4cl9dY
KimnMdms6Um1M0Njg/s5pOXinXaP2VUkjNb03uWZDCEVUV/P9xTxgYwGNJJq8EEbNDUI6Zg8dXaZ
+iIIAS+9l6M1EHH+JnsrDI66deSGgBV2/CuAcd/iwLPaKW327iORg7S1mgCb5yADQuCsSu2w9vya
8k6kzcl1aN8IsUTGJBY7YM9BDEzJLXATB0r3sD40ENOo0H4mbIuXqC9Ll0L7q9u0xEF5B4X3IxsE
lg0gK291E/I73QjKn2VLBF2eWUndHttpnFi55yvs3FPQW+miQNFmKi9hNH1S6uZ3Avr1aoUaXrUn
/Qz4n8Y9R0yGro6ZwcZ8eM1EHQmtlfI0QB9kM8Kwodh3ryAEoCep+eFNb3Sl7tW+Uxx8Gqav8bwW
zKJRPUjP+dO3fUQpDfzHx0s1WAR0Ph0TCTV8l0PlbON+chhYG5XUjcMnjhLR/svn7hB65UHp2V+b
3ED5KnkhSf09pntfVcYAcHa7N7/xoRMJyE8LxDdTBhDy8FDD+3meJgCs1y1X/zGooeF8uB/QEgnG
xI1ZlcjZsGWIHpcgkI2KLEq/BTW6MN1qzJyRxbmRWE4DgEcFmFaDdF8j0G1EoDW4T6884+J/vCE9
rGnDzUPTarsT0z+78XlQayxa1VNxLbAUmy/p2+o53FoIqxn05QPD/XM0FCXJr6FBosOmzUc8uErH
gNt9NatmHP9n1KhjcrRL/B8vuEgTqLtI2oxKgs17UQSJlkBf9L2rdl1mAkz0wcHk8+G8r5MvHzRS
AalGvxvChzGqZVVp5tV2TPh2t194bWgYepQ9wFDMtv7qsdrA+9nE7832p7Zo2iAJ2sc9vn7eTwW0
CIecsveub6tAvuqkpQ+eDMxImu4z3U3dWf1JDGo3HDEspq+jSBSiFBkhvRvfcQcyqwt8aOsGfx8m
8wKGgoNN5a5CUjT0xAUk7YHQ3EcvVNSix7Wqlowb+Uyet5uXuqdG5lnsaj2P2OETyJW3kbFDIcT4
ak969ZJq9OscI8GtvbNRLfNsaVY7nfxnC3wY4fQnxuQfjp+p4YqCB14ifU4pbPRUMN03ENWHPIxJ
7xOS2cZh1/q6YSvWe7tN9Uy3Enx/rzAdOV/vd2Ui16v7KtTZJ0J0c5kIMqGt8Mmbl/sI4NOCSnOa
1+39s3Y/8qx1FUugHOsRhxoH3m9FGhEIdHr3nodRpNEAbLm2c3InRNZzG0RaqZLOXPYafRXkWf3Z
FLsqWxZU+Yy4iMflbX6wWcJaOcAgqxhAJ3ObdduZ8gngeNl39jjb9GIg0O9HGeKdmqy0VVj/Nb1O
Hs656S0bCtuR4dND/bSxvLQZoVX7QxekhmmyFVPFGPd/Lpq+ow2PKLm69Cojec7P0RDEXHurkR45
0ZQ9Ka570NjILmrQRpWSPiFv3yyRS6DLesjSI0f/DT1mkhbPk7C8GPbJ3dGbFGN0xQJVrKS9Y0/d
brbru9g7wjls23I8lfTkdFMhdXE8jDHDUBVzSz2sQ/UMNYOta38rUgVRBjkJv8CJ2i+I/5XX9l16
oveeiZBqe39snGuGJCpjm67/3ereWXfhwElgbChpA6NjgZ8AdycqsiyQmgG6KDVzBP9jKWVJwWrm
PGw+qRZmjiHzMV+JX8AvsQvl3Rkto28Kc0M1bynzlX6+u+D3pOTGC9Ipm4GnxcQcJSWk+OQFklqs
nt0JAyFp5RxgV4VX+jtMclTeqw13Lbw52U4mehFaE5RRovFWqFpjhiMo3uLsWKoTehrw+PcAjl8x
xt5UVs21rXlMv9r7G6uMNslLAFJNcLf3s6CB2KMJYVz9V4M4xtplZ+lwWUy9snNa3RRc5APhGX8U
bEjYEjcxMpXv6X5NbxSco+eJHXmjiE6tkKtgA0EGg7aQxWzsdZhVEoseFzM2oxWGsF9sozY0v5TD
yDMZmTuBX1LLgFbFbp31dGoGEJrK12rY44BjcX2xafduG/VBBHpqwZ/MgPEDxHuNYU53lsUt8FRt
99FoqTN1+zSxflT0KXqNHwwZ7dVYwfDQc8+ZNNSbt0wEhrz9BPeDqDZ69+ov/OBA5qv5HLj2FA0t
HQceZtNSy9QC7oEyyFiaOX+Dd3AXnZosHTWQxiy7Fcu+PQ1wETO8Jdmn12QY6hnVXdmevXA6gEXz
8QXF/uGc99HvkGnjTVQo78lF2gFd0DW+ZCHtgWEAkmkWpvK1OylPxhzPLGees65E0Kc/BCkT5WBS
fpkVhUNSoVvKkOikQxoPtYWYk7mwdqEry5Bdfjit6yllNfCy/kisMm56DyTLJv7/gJc/vdD3iVXV
HNfK+D9TQBxqHwAhPbNObeJ2PfO+EM8KdwjYPb+mh1za8eLaT3Q3XShpCL7FIBYoPt6bb2I3gHtq
RrbZYN91m+UYZSvloL806oJVmshOI5s4xPH9Q13wZx7HbNlJ+elwFJQFDdIin8cXTSigZhICXOmi
boPYeHk2jLLspqtDRolyNXpH50vNM4NR7Dk7P26pBkxFHn0QEK5QvdFuBiQ4QlNsFCGZdDRPqllk
gLPa2O/JkPws/JdYMVdLg1Ksc39vzPNaZVbZT6VjsTHEmjquQY+Aly5ccI1FZvvsaJRPSMtUtYYS
gYbs9GNZYUwnww2BWN/ORJBGliq+5MAFtI1gOjEezn8qGL1eSw4lXNqUgUSQEtVCd1TUlyUGCx9h
S4bYl9YoaDniXHgX9V12Ama9gQJnbYOWZUfQRPy1fMF/QqIv9M5ROC0TCrOP0TKbGOFy2kil6TaT
MP0GL1RsaC+x43tDRF1lwkpZnmlLXbIGIL9O5JM3yQMhYny6pP9Iny5CIe5jwNzwxjb8qDlPsyXZ
LrgYK3Wrcu0SjNA2IaVjSNdgZ1yDQ1wnAc6m+3qV24gILpctFRImYGfFOCbg2Jme8OIy/+zxpNtD
oQwJg+U9gK5wSYrANS0HzpgN6nFCcXZ2pRUdZykuWrebDo/hWNev3HM9kbKKDkYgAUrPbEUNCh8a
kQGjeRf362nb5+ZvkqEeT+Vi7d7EkIIUqxJjpr7ykPHbqPUwXeRKHzvwBIXqzy9QVYCz2QoUqeye
OWNtLRkBaTOF06Cu3QUQGF2LvRZvu5aqZI962mOF73GQFaOsI6K2M+n4TnxDP9dheuQJtNW469nn
pCMIR12lfH1RGiH5dVK8aKTmqAbAv+0wOlGZ71c+iW9mxaCpw9m58wvFuqVeEt6YKNIfwD/1/thX
WPRgTGzXjaUE6YuHIdea4kO94gX1awHzP/7Ezg2TGUpcf0WWppdNCXHyGuwMjsOg8VfEBgvx+mY+
FTyRR6P0ABz0F+uSHru6KwI6YMAWTfSqoU2nwNHOA9k6XWTvAhuB8UMFkN0cL5Rb9bhX8JZc4aiW
IyjqNLGL3wo6d8qxtjcqlv1pIA7Cb7vVDjPsvKx2X3fEcQXAWFkcVCITMihQXlszGviIQ8bMXAJJ
9rsNGdJG8+7oxFf+u7htnTOe0SBUbrBeIsVN3EAE3ZPKIaBDOCCnYBd2ZRoiyCXQf4sxrWc5uvF0
23yXOKP8YR9f1S2bjSXaHmxKU+WFH32jiICAV57YTimE0vEuRkNF2/W8uuGp5wyD+ZWnReaRZFu7
gLHe9z3f1BOiZSUjIxyUKk0nMykVeVDB7/DMcKfkixDkkdA0eOn6RweE0sgnLrSAQB09ofgimbBY
JRIDibtFH4/GsWVk9Jj+VFaTMHni2Qp78gmS+GTwIp1qA4bSKdIoe3wTpo5Fi62eGNsiQb7tVdYP
fjxj9DUG4/7tl0/OtRtFyEnd7gF6JS0KC91Otd+tegjKr4OaMAKDZjGo36s0iJ3nEJkwb165n6R5
yFPzg5A0vBHBoLFWS6RCHml14ztSiUKH8QDSZjeEle+ZEuwm3DCQ7VGSBeFcj+pf9FldHSVc2duO
a1XwzD2G3jjlWAibIQZpqLIHJXtMA4CbRU8Ym4lAluSyF1QitgcRM25+be7R5N+wq57SHeH9Guq1
cxiWmvNhsr188jfUXpt61WTj6E1c+lfkWXpIKQG/MxZbqs/IwzURGsR0WwKozGihsLIu8Aba8vLs
YZbZDgH6QdFN+2FJ8/ztF8NuMEzZEAVvXMhwJFLVwYVgTe/YoKyw2OKnKe1z7LsZEFGBTPjKiUC5
sGF10DTYK/Ej3woHP8sPGhoacDlVTqqoJJ4OVE8SQEkIjQKSak0ktgnU35JpDJDwyzUpQQl0K8AB
ewacFooJNQQaVZ2U0hfdPxdnREiMMbp+lW9q1jDDNIfQol9y11p4FiKXCxABmGmzKK+DNhNfr0jz
FA9EayDvpUcYsrLWykYR2tKzDZt5SMY2gO7wB4hEzQusfUXdlBuSzlIYLwnemJAJjJPippcOATFu
cpPcscGSAbJc20jYpqByxzqnN8ePpqaWddkg1XNo0halfNzKlOHcAnq/gaQDwq3Nt3twQd5vrEB5
2TMdWUkNXeLNlTCgl/QqMzYKbKzdTXH0qY4DHqpiSZM6HiKDur4BZ2upmkJyvILuwvpwk9TM2ibj
57TG7GLdbEcZq/B/AJRbmam+gOk0EWeWWXdB4uPGOuaXSF3lYDtVee21y29+c41CpefrY7fNgPaO
vhFE8VsYnkAqiDK+OgWfExZEEHDvFJSX6PQdgI0/hgVMUZ97ETI/xk+5VPhu9Y95BVFuNXa4SwGg
bn4c0fRseT5kecPqIVBzPxoXok2vhl8EdGDZnlwheLoxYERlBG065nUHCKcjZuuUTuIuHEKeXZQU
b+HGIVGnHvOcOr6bGQfl4VMss2YQnINcxJLPKSfF7ZtX4+1/Ihnfh5Vuf1/hqjAwCIDzEPkv1ygL
nKJhNjsuhleEhCM6DLxyFRtmTMp2423MVzjYPhGa59dGDXnDw44Xw2dIomKKadMVuTBqAGGq+zX5
7YYpFdtl2Nnwn1hmFevNspx9GDNTCQkWriMFphOefV1vnz6n+KoibvBtIKc8KDa/+7pHiMil2VUL
HD3ueWnUjWyLhjn23y5ZaaoOiXSNI86BEaUokVqL2tDJSjqFnBZNwJNddbuvuRiN7U1ShkurcKJw
KD/z8rT2Exy7WE/ajDfyxrt+DvGrjQB/PKfK3ACGWDcZ4s1Jw9IC/gb+OZ7WkV3wp0A9v+j3jJnx
juCI1DhQsiAMkOe0ubds1QigLzJo1AQQ0Gs+ZLtwelYl0Qvw34xQJK5veXsp0OlkPxYDxhhZx1Pj
6vP+RbOeLG4AmdTVKkoDVTUlknsl7OBSJt0OYiNwtz8dZxw1AP7tZWSzr7/O3JZqrrWL5DJSlRje
N5LODrQVl438tvyZUJGOZQAwR+7lhFh0i3IecGlaz5IvCFGAAv/h4wqX6BBr+bkR3Q04ljqU8oxA
9pb3H4r5VYpBFW+A4AD3Baiyzcqf37TeP60c+NFkPZZai/kz4edkqCnT79UkcaYNw6hGyKiYxHtC
aJ6GMPXbrdp74t0N1P5cP12dX76IsgVgp2IdJCCzYZjAmchl5vtyR8o1/ViE+eyokYcHRu6k65Nn
ySCNiDeFohIiKtpi355NajSffZlKiuT9eTUQPgcwMr80hsZ9cCsYmCChX6WNsuO5YltemlcQmTBv
35M9/nKsjTmRwau/THf22q9IXZKtsmA0wEsJyX4EkcZEYe32UTERuRDof1JY0NlTUj0vVPcsfJbU
garv7APvFB8WiSnD5BqOrfuKr7iAeDCJN4pd4jk39F7KmglWHFSukE7CLSKGKBxXApDwLU8Yt7B9
0ZefqODHDqMd7hoh+3uKMoMWlO57jyTv0dO4aZPrK1Byo+qESYQybOMU/oLLjx2Ir8ZgF7X5F3Ie
YusAN/sJPoUesHIMW6uYTycUtoVqaBXkstBcN2ooAc5QOaTJNmNOhxkN7bceQGu7UheJM9z1sqPH
6kwRDhpjNzIcxiXKN8TS3HNvxOsjiHWShBXVE0GjIrm5ldWjmeEr792Q1OOb58bbD3yLkgAYdmc+
FX2whYKh3SvuH1e8t+JzVR80Q0Nva0K9AKXNgmBgsCN8ST6t5GxE+grjZE8cMB1Gq9lSSWT+LgK7
hj6Pm29YwDca4DSwA1q6sZn+FZwcHq150HIQcUz/fCiFoDfH8UA1sTGpP1VJcuRcPYZvnCy8JLw3
u61Vxako9HokPQXUT8i4W4BfyRIgrbJrNI26LL3aC3mnbb2VF53ZNNwd6UCx3Q3RlVW/7JD9G9Ls
Y+gH3r4bdAC93cRd/bokmvCrUITBoXdg3JD/uryteukH8e6KgifPrxqEKG/M50Ew29oNBUnGBiEK
wa76FAFMOdP3BVxNugz8u7u+tw4L5BAXavhKX4CKEafbUg67IdippM7qzIPETz3XS32CVhj2KI5e
K9gM3SDWjyYi1Cmd/6j/daRfFwPXGAeq9nbwElAac3m9UYrFDSX+7IA5ogcvuwM3FVzO1bX6qGcZ
xnENcPKj8THor4o2wkW537NI3r3F6m+0zZG786zg++ImEI1QzGVr8WGV2Rt5erKC3BqTIyol9Ad9
4v7tpIU6NdaenybWQNVoGIy9oPYnklI0oulW9W2NR5c8LT6880TMB0wGQQx2rqbG/lC/7hMBWu/0
JY7yCI5sh87hNdFSr4asra2R4dupjlXcGqh9lddgs4pAK1dt0d/pZfnxZPWfg6nY4xRRVe6A33og
2LBPD8FrrAQFJWB2/MzXfqgu8/28E3CJNnXURleAsFNgOQ6Jjf+jxOX0o5MsfdELZjXK+DxkjOv3
6xtmqJP1rV/FDCXqWI8EnoU+lAJqhnXpWARJE3lR+l0z7+IKNfdkyZ6lGnZFf05Xim8PQWRPbq2S
d3NheHtmezhfu2yd9CmC8YRg6GJG50bpoId7FnJH7VoNL+Fchx4cqrTQLcuTTGEXNA9NMBfqgrPV
rFxe7A7Tam6j/n5BaOrpW+l5pkvYYUp4BdHau/rhhHeQEhnVTzZ9eWuII8KQlTcwOaF8wfVDs73O
wYkElLhbEWrgaHycRy8Fh784FVSPrOISmeiLf6Uc2GLYVC4AivGCHgkWsfW5b8Pb711mpJnwbDWI
CnekTeRY1rsY3/fS4E473XnUl/L6lLGjuxJ6d8eRfYpH6TtDGr8OwRIOro47hbu7ETAFXkrggHx2
xT6sTjNltO88hT/3g9VMqwaK8fMgMCXww8mSDquqZS1I4OgYQecGRnF5zVFgYSIz6GuT3Vo487ar
NyBJ/GsscBbffVxmpYqGc04pNlNbQRVORJEM7gSZMXhtTIupG863VIooxLMMLB500EmigdYipQea
18UZGyymY8ZSSET5fxnPibjkmuFnxk9nv+FaiVLYmQpXYKShpvgRdPK4jZMgFWIziRvU/1DhBYqy
hVyrBQDDhTh2wiDNi2VbYhC+t7b2j+C37jPXDoYYQMW+j5dufweeC9BDsTYv2U0irsyDlorbJx/w
ePFAw0SK7xgnn0tjvDVoCkaqWIz2CFwsmXpnS4ryekxTNPSUJl+Cq8yEO/Q8HBCxIwaAj52dBs0X
LkyjezDcUhFIuYMKZTc645UXV0nSlGJ8XPtALOFCYcxsziO35klsEjKPEs/LtGmWDdiW6+GbK12A
WGV4ncFbcdylOs1H1nTdmi1zeAvr5TDIKXMJv59iEb/tc+23YoyuFT7/FQzaDIiSHYFfBzxt6EqX
/xbAY0sFKRtUAKE9A4sUlHND++yMV5eDcOiDiwJrUt6MBHe+4qHMVqML8BKS0oVFveHHOItFrf2u
CF33HXpC1viX9NKUbpwi1aFFEu8vwxkxEQyLhcreuvO1afELdHecuhKxRMCUmv9F9yLZsjsa4nbI
0RZpdpDKeem5OY22/K1W/FVLPnhZ1xiLj7H9Yqi5uiQwqKGky84PidA2/bKTq/QD45nPz9ioAvja
TBYVyxhyR3HDJLMRnkUEaAhozG0T9dH2ayysYqT2OFwmTfI4krf8+vFjKZBVeRdOw13K2RAN0k0B
f+8PecaHubhnjKmkN+fzeHslplr2qhWkAzkcsMB9WIC024N22/FgW+i0Y4xFBdUaHEZQ+V8VATpe
Ui5v4tB2uO8H5p4aJJpbOC1Ob3NDamjgBcahY+Z1/VFuJtLl4/gv1DU06pPMuigRyps1zmhETddC
qhFKA9HxRz566fvUdY6yX+xNFAEkFZ5riPPYeBv47StTnQObPH0+lv4GSKtNznFI0Sqzz2oDFkG/
JtIHghF8g4nC1vYRWx24X03TROJnSYUO9QKgjaAInVcVBhCF2krRmvGAauHKZfWipS6+Si3MO8KO
duKR1jibaKKY5a6Llvhkb9JjwMwZECsqrj4C8vgIvYyluqrGL3EV2Er9/SSWzYt4FHpzJxAWdZ2o
DkKaPbWE57zOXr1XvgpsFQv1Z1j/TNtfU9ac1muPDygC8dXFNOZ5UQtBCfho/qj6Bj0D9refcrTh
4kxeJtg2kDiPps2SmFTqTG0aGCbToAWqKGl8SukzVwNXB9KJCgCYHRV9FzuA2PHTQHHVsU+e2Tfi
ICM3LVmuQYWdoS7km1+iDibC3wavs/HzQTbsiz/dZLABjbMbAW0gMfU0cH1wPWbPnCG8sKiTdrFd
kOu182Ys4XLiRfqFacjqAXMZF2ej5T6jC0qVvFdY/UYfhIBy0GwjOZAewGI8GvaKVv5lchcCFgVd
W6uM9xae+QDHydKF79cK84q4dnPpiJRnGj4WVYexPncEK0J/jtp46ox9UT1q3BHSzrU8pAAOCb7h
JbdWObwBCLOFTUd+z/aRwaZ7IVoyYF/X7JS1kHqIXVAP2NlWyy7212OtpB60XfHHMvZ3RH6iGKns
K2KNEjhFo9AmEcMUqVL1BGJnr8T401GKtZMNy3PVQ6JL2Un/WlpoI+fpFkTRomrHqDe2+qJdb/1O
pgRf20maoVmNVfQx8a5GKSwmHLyEDtV+joyEQPyflLu3GkWUFU8mrEdMjPXok+jjJwOtUE25eZSh
PNd7XQlaLPC2yLUjWEMYNP9xP/b60y95jdXkJhzVwD2SAiIOhiIl8GGYRkBsMcEZaelVNE7qhA+r
svU0y8Rz/YC3HaoazYsRPWh/ljcFIlaQhVnonoiDRsNAfPttDB4bJMbrJTSD+7UoelJVv4wwrIV5
0Wr0nK34+gbL+qMSqqk0qneYmeHENnAQUDHvUFf5wORDvI/VsO6LGbZdDqnvEY5Wth42vR9K+0ok
5VMITfvtNe6CC/heRUEKlBMak9EC2iNXX5J8HsecJaaqOairU4KiHE5fyFqjZ8Q+kO8vL8nureAf
Xb0bZatUCWd9a55MtJrAm5waOty2QQONj4RY8PG2g5ipFni/T6hw8itA/gdK/cTTrcW3Z+R26KI8
m9UHDU/XiQmmRSVm4nhna/rH5o5io9Vggh7ms31Y42FtOE8zGtfvjTm5ZrbjJKEoJ5ch2ZmQR1CR
4HxE18DdGAUHIVji2B+vYs2eCUVyvG2lQ49uYDq8lzBbarMeMXAA7tqQ3Ev5EsdTu0Go1VGF9PUY
NsyiaLfGGvsnIP9YU6WZUVTpZIl9BORtH+JObYLjWr0RIbBPMrfBjzbQuuwE2FrPpyYRurLLyWqq
m6nWEmrs3aIvSh3Rz7eK9baxz+NuuHUKiuooMgcBIKFBysUA1El4t876+hNOqZIxzqMG/A8cpdVh
sq8r3oCtY0i6hNt1Cd3nfzWUYlWZSqEOsWxoxOU0/UpDm5C40OlA9UoZB7zgx0JyOyNYnrjcliYw
FVk/6MS7sYi8ZGyDAlWNeYD/Jwbdg2mqeUgnWcazIL409qJ47VpRTbg3et+k5mZ/+3p7IyHj+gfR
QnXPgD65RwTcMAcOAm2ZWVPWRwJLmwxuYoNcASHjavwtr1qkT+q0mbmcKDUWhNOT/oNHMpP1BSmW
dSaLS7pny4ZzVdi4/2QZ64Zh9eQiZ4xQRx1hQCZUf1YdqHUZHmrmOESnw8zto8xNqFBTQxeoZ4Qi
k9uic4cRNtbF4wB83GVtKyhmvEdMHsq0rZ/O6OowjM8agJrak7lSEUxevO7LbubkJuEg/ofhMENm
u81HKAMmrq1E5YX7v0N0+rzBXnurkb+IhGOt3ObPljHuP/leOvzV3ifBBgm7
`protect end_protected
