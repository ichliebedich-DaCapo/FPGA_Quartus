-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wmHGoRtFjXKUmyfyszQvuBGIOnH3LBSe6eJbXBvdUcGe7dZBgFRQ+4lngAmX2LPEeMps8by6MPv0
MWpBZ7lulsCzr2a7rjAbczQfCAQRiouH25a9PaOGuyVlbVsKdA+ktfsfbXof4d96xOyOzGY3zkG9
FkaK5rFVJ2oEBMqU4HQqtxx0R7hrwN7zzcTYVirYcJkHaz2PH5CMUWzgRlkhmFsqx7ft+pRLQRlM
uMnd6XTGjQF7IZccK9ZGmKlVhY3XcrSLY0bHdRFzrI8lVu0sFlnTAqvcTDE5PiCNm4RqNcwkGu84
XQeel0IHY3ilf+6w90JgpR/sXEUs6X7uhD4DvQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7808)
`protect data_block
y5+wb56mQrkoj07TJ8aY3e58dM8iJR+OojrQv7BWyNOE2mIOEX8JwRza3HcGUoLf0JBX6AHiZTUR
kmHTD2LZS+jFIpRMvDTfRy+K9iyD49iXSPRuOhSgth7yAw8AVnzU9ZZNdstp8N6ixaH4SoNihYVT
DRRxspOdUAYxBIv+lCyxCWEM9WXjd5GrcnXs6NlPtXv9cbejdXbrLLfKt3ro94lZgx6jkT9d2qMo
X2FfjZTVnXbgtBJAtuahNK+Sc56VKqPxptECWKi0X7PQSIfde3anOZNXoYVt9y9CumDek3xnKEoc
NiIs1nyYbvOtM5eEhx6hesRqDSZaR8yXPotKsQNv9mgMuPZ1SPLQA0mvKkfHih+Oy0zJKj5X6CtM
kDiBsYPjLKoXhracLhGMyG/4JEWj7h8dtnSmJUWV0egfAuUDTOCYldlZQAkhaJk13Q859Cyreqe1
J69C7fuD+4emfbUaRaCY+EaGjeUzy+ILQR89NaULyl2JfbJClOjsfAfat74/d4dX2n64Uw9HQIGv
omHlkIZjIcIVvuORPqsSowkQp9FCIaXonCL8yxAOEjomX0NMFi3pRXQF1wT+K1XtaBgSkm48z1Kj
AvZFKS2n5YvctEpQML4H7ZOZPs8Fbsm4/fxtldS+Hwkoz5acN2+/sJrhjtZZfxxGAD6FzLbNdHpn
2lGIPtIQDX/Ao22AQW6PxvNeLjhfJPOK6dkbBC50o6fEwOuQnBwCb0n/YP4Q4ZVYqVlwvjTSMUCO
IRolo5UPZSWsCpnIld/i6s8DNeQrA+zC29U1p317oqPqwfET0TQZcVN0d0hHAfSQJdbR+Ub4+vAa
bxe3a4oI5QwRS3f12dRi2w04N7k4R7XMyxC96WM3NGH8nQlENbwUxjVLz0l0onsTriIPM1X1ZqaB
FRfdatVD54GQLhsbroldeLU9sbbqzvmBBGdbY/RDHdkDoYT2ii+/cTjusrlVAWQnPTYMzv3Y8wjF
74pdvFpdXgbkZlcpRUBYy/CThj/Fyso973PhKAnKu4EXfnwEgn77tf6v6h4G8PmFQiOu4Yq55e0b
g7wf+50MAkNQKnhe23AzB4fhkWdyWfIQtRNLGINRVTvwffgh2dinjB91atC34a3RDGnw/wzEUKO2
M56vEvjaei308QpssdiR6Fi8GlBuNtnQWAxWhFGSUUa8bqNX8VP2FbjruYDrQ61GdACU8atglsSP
ie0QboCPPJQFmx5X46yptxkes/qEmj3IeYcJSLiI247KIYcipmYQg65PwKPjzotVDHId2fqzzzc+
kmkaR/QN5plWEzuNCaSpQjliOAS9xmFk0rBNQ/B3emJ/m0j2lFPDCriYMpMcfqjm+okvBcZ6sGLy
e/0l3GauKuX5PW/WO7TmF6NZkXTbT3rHHlijPYgsGRRiwRr4E4L0gMVicBZiDaP1KMBS9YwZ2Zn4
NinudhM05/CULVzyVzYpsbT9aN3FiIAnJiLY8GFUzo4qP66nmYJFX7jpuKMAUsaEETbFcL6nRmW+
MzgqMXH3BfzBRWXObdiyuWx+5FVdsnKMNhZn4T+yfCLbBid6wsx+0up5eHXLeSUurqWC7r9wy5Y3
hXiWsPEfKq6sMVuhH54+VsW/WJyjk9W7aDMylpUDR7Pq/08gBc9rdBCVMhOmM/BoVDHwVOf+TGtA
1ON7bzO+v1Cd9lYMKRtasZGnuthhZhIKC+KIcngnTbirIGn02jl252tmhZ7fv603TVRq5T1guj87
YPXuGK6YTsx3bbODigJrTgm6EUjWJ2x9b262ve/MnJ9t64Lw6axmL1rdlYGKxi3HxOveCv5e8kQi
EKmnxt3kyuzZL0bUnwNI3Wt30QuBys29V44ghYYYnu7ozB3B065Z3+MQHQpBfHyP9pbuhJjWIixd
B/X35h4BBa0083+akYH4nyYrsVRlcIPxeBzrmLPcaC4AR+29doA3TNsUeFf8G42Wszt/iOyN+p5N
aYoIstkk38ZVKRR5zZMtnEqZNkohdntlbiNz6BnsEt07kO4v1LU3/jg9f7hjXvXTbGnIiIuyxbV6
JB7YP5i280VmJIBdV39Y2J0PCQEnUL3XoAgZfxmEkujk478UQNlqpVW4NMlPxLoloyCnzSUYlW8w
e4KltHSGGrQ2v2ARwgmScMdZiJU8YdbKSMiMCj7slpZ/w7pzRyi6N4OFNa4ZU0KZ4i8wwQGOTEoi
gF26QpGf4ckSpIsTstpKOwwJuYwE+YdOHFLFtiV+LtmEbGpSQTQMOy+XLU1Ohl3ig6hQDs0Io5jO
jbD3XmAu5km5P54wL21juTp4hEMYz1Z+2ON/z7qZHSUGTTQ32JMRoiPXgfIlt7KtcuI0GF58rbxe
Pfvgci/B9vCniUgwxFp3I64iKNwljY5Mp/mjVsJ1OtmOIjNvCXY08pKHPcniW0X3Ga5vZI8fv07i
bEshMjTp82kXyF/SNGGCkpB1cndmSKxzmNeQoj5FVZIgMEnq12CJr4SFcbjkygYsiaYbZsjp+nEv
yMo0xyxPuwlp0FbNOt3jZ52Yy7QmI0lXcJNZDvSIopCCH1MWw9G1NMAn2nPg0mQQDkM+NGYJbCUm
abzsqN+xf+wzO3NGcmcay/+6W9d2bI2Fb1D33Kbx/Y/48EVTo6MWaHPDUxpDEC65pJ0J/W47mv2n
3ouXz46t/zptsg8C7hHi9+NCdLsbVEBhe1tR5DQvSDXS2Pu22s7Yy4jVCKqn76ykpmEwUN6Ial+t
5pUdUjG6CG4bMCz2ibWZLoLf/RFLJf4wOKuGqrZwKexpqbI49/D2/nBXPgPaPyEodzAdYt7jG66A
kLDD6vvr9BRAQq4ZML50JxL/ktN9Zjid1vY1oMdwiOLrlOEInyACebNJ1o0YlsAMWz7G+vk3HFrQ
O/LYYvs88bBXxgWgUrQNPpTUhgusS2tnEN/4FVKKVd9LpuzF1qUjm0DksnIefTCrdE02SQt+oqIl
eVwa3X/OejGIhQwiQEroUfOuN1d1VgOaH0UxB0PUI8f73gZhj8jMITyGM/64+caqc1KlfmR3g1Ih
cm7u4vbwrGmmAzd7UlqQFc6Oy0Az/tqIqRf46NKQlHUhbFoCYSu44hRLHVVZpiQ7kwsl0mdDOpD0
DxlX/zjqlRK6lICMPwJxm1NvlSelKmUwfWzeHQkmLt0Hxsap97mVkBJ+Un0ecMj39P7JqxeCzBWT
uHnehvaB3B+LQAO5JqlI8X6AfkZfjYDTpPMOfKwK6oPNwmzS4y5WRoc3Vi5+Hccg06P73+cOUoq3
WNMz4/TTWNzLV0XVeOBeXwzd2SU+YDvA+0H7n36g8thWBgptAGZnfDza1Uew0bYZ2znCjfSZGm5u
Vr2i3Y9pckOY4ENYjAIVeE84FpIHMxuvjn3vPAd7BZb9k9aLXzVRokko2rwayNZgjP1se+Qi9ze5
EJmCNRmRA5iytVq7fhFZZpzIzxIlqbpUWFaKYH0S/FgBnr3FdN45hSuZWYgJRaGHrUpxhheWfZL6
xD1B6RuT1btaZuC22YFA+1sB0GWOO0dofsFCySZx8o/MBBRCrTxd7uY/9aVG/1CUsZD0RnsJMU+/
duPmW4nLsKch/2cDcQsX4mWK41Hsm4Mo41ZtN6C6+FQgPR38YWVDP/MPn+gySSHdeMQSLuOwRB+j
am2cEPMrMnBPnDdbzJrJzupl7GarOFZwf0SLiJyRQ2Qm2swQ4T3nIE8YOjeVX1GBVrA15VF3lDnh
4dFtf6VoEHHbK4jiKM2AreGvccLa4Bvr96H60mJS3fPCZKUYaw6esLDkK0JEKpX7nFOenCNepEK+
NCAxZEOi8FApvWwtNTOyhQ4GyAABu9kAiALrTji0xCl2p7siD+Uup49/+8xMz3uFcMkRvVygdBlQ
VqCQk08UfydHRYSfwkuPJUqr17kWl3YHcqGnLO++toVMqg0sxnAiXrMUfx6YKiVWfmRxK4L7EgMj
dZJX8P2eoxMNobXilMzLKANelCaetjK5Nn2SiYSgcvsa8wRvuW3qWe9xiErJVxJj+5PL1UWr4QzS
2i3HA5en7iaszlCUPQtsepYdE3gFWMCnjdBgzgHS1ZJYedJ0KZkYc92FWzHwSHH9h1IGc2KNFRde
vqnMlwFlEp/hb7ssjEAm2ASxKXaMsxRSujG11PvO9Q/WdCuTf3t1PKVKloqHwO3JtLOgaBq9ns2e
t74gRc5OCmQ2aTfqDg+s0fjT82Ou+pph/XeRmzRupAAudGR4LR74Fhp4r0MXUbjsfaadhx22LSGr
eCfZYzkgrX4UN/kqZ6pOFoAxz1wwRL8gHlpZonD9FmTc8mq0VUaMjCe7t7CckE9ZVwT2xlMD6Nfu
JDd47turrPX6dI2yTUW6j/CzRYPwNqLl28sT/k1sn0AsEl3Oa4CgXQH6ttZtejOYe7LwdBFrS8It
7qR/BaRHN2VfMXOwUPkCCImxUHhIb5bYUEB/WKZSzqUJHQCxmR9cAeX00zeRm/ECfXDwHIRNiaJh
czx57VaK1CWftfYuY7m9TOAJxFOLDSuOlet3z3WxR7wFu5R8t73SN/jbcKuZdnLNUv28HA0VYByb
bJuPtZOD5qLSzUD//cXTixFNk+YFiNhe28DO4Iwmx76YckLw6ajkeW0lSUMwKGVmrUWIAbrLBf+n
uyqD1U7rWOTO4z8/UTiRifdxmxELoigi1lrYtO2jA8sruje6htD4XXRyIz0Ruvj4MJQ3/1jWyzov
1ABVbKICnQRDyfZ1+sSuMdC1PDkyPLthtVa6P3qOFMd9AZzmuEKcF6YaKmLB7tbkE1gkDrR0jpgr
2gTjKDE5xSM8nT7ZTiCkVA4L6DedrNdWyLM6LsSXq8VylYxWX5dtxa69Yy+eJ3iQN3OlaRPIoT24
cQOufnQenlmKWh5sqgC4ZGnK5M3sYtBNNqTjm9ZNJkG0HFRmfaTa1VLPYaU0I5Pbxvdvh5uEFAhU
5f41GZouPd/tUVZTfoRV/nvQ9nCDkgTPjgU671WanJ1uleiI6RGZyzEag/yF7L9F8G1IXacNuIdn
DYsHZpJJ6q6jdurWYE0CsWW2/LBRk2yWnEw7kxP0QQLEQpdX0czNAGu6iZfwyUZF7ZcTTuYVe+PX
vQVcGnvgU2ZTpA4iPMzTalGfgL+84OuDSUmUtxbz5P7J2O2W7jYSPCP4eiC2DWpkG1gc/Zca3fF7
8ni4uh1+HO6/lp7Bgv0nTYoa+5GX1ME0Nz1/nbNve1Ml732YV6ugKzEVOIsQw2KWig74Cgv3J35n
fxCg+vxjqN7rSp6SQbs19v24cS06uwz3pVGCj7OdlM9Q2MoQSAurgqYbOUYpbuLJIlwbj7aECUaO
4Dvm8pRhkOTehMRSKVNlOXj8Xzkz1c1Q/iFo2tD59oLXQmq6QQbDzbxKJsDoZAPgg5EA2a2Y/nBs
2I2E7zbNnV6JC5Bb6RfFa47FPA+qMTO3NGSK2QUlXyEopPs83bCSLstKkFVbri2mR7v981VUnqML
OdicArBPWhaxjeAjYYIAzNKstO9+VWST7WSWIs+HrmgKpYyV8r7yxh+06tkqOKdsJE5ftbmu6oBJ
KpwkH4V50jV+jmd8CXm/18+C57Mco/xc72EqJgeB9pRqLlzuMwU332nbZgaHsqw0msEuz+/8SmRc
UTts9S+o7bDO69nHRHLuwhl3KJ9yFHSw3t4qfneqR3sCJuKyRvyfvPeYZuUtt6q/Zp2zkJmH2I+h
kqr8U5zm16liZh8ygZmSmvPRzfHy/3Z+Ma6+kxk1IyAxJ161JRav0lLh2H0ccjsZ1qnLs1X8zoSD
5HbbhPryQpCRRuko3Z3uuilbi6kw7iyOFHly+FOgdcE9TLjpRQ5BMsYh/uoA92YYmkAKgyBoTewT
3XpWURRpgKRp9NFOUOrZzqgqFK5KiF0fdwah2W0/++TvD+O/olX1XX8sTj1UQo1KLXcebymeoBIb
14Hp6IW/wePLnc7Dqqv6+R67YLcCMhwVqNBIaX0O35u4liTw3ypb4RlIrKA2Dfmg+LbGWAhyuib0
S3wnCHPsncxrhQKEKW3vBcrC/aOijKhG8hUAHQ2eJ6z+9cjct1kwREYD/fB+/sAnBFtOZaF/WCwy
ZCsHH/5ZrQ6FI8PjxYG8qjn8LsUdBYF64Xso/6cwqamIKGBMdgXhpvRwUtRJNnP9+yHMTZ1mgrvQ
Z5dBWSnv3M4sbr2Q31fQdVH+PHNwQq+3G0sFMNXZiLfXGRBMKLRh3nexbc8h1HF2y9KX7jkNKsfT
8+SMQlwPQEzoL3O3mLniR9RQBwKrsOsoFr+2V8m9x96r2KUbgUc7EeBVlaqv4R4dUVa5Ac5hkXV9
qgfOe1Z3Kb9jDZioevXXGxgErprw0kg5BboSCHXPmgc6MLiH1W4Ra9iIE2OT05N4j1ChDi+ZAW4z
CFhB1EQKZwDZBeIPYn0ypogdaAlQbL7Mor25me2mWEOoPu5JkYXlpDiZO48d1/Eagy9943gKfTAt
scNjdXUAb5LzNI9ZLSMJhq3CS1x1ZkX3LZbVKX615qbJSWIvngkDZWN55W8aXyoQUwynZg/zuHRw
Z5JNp+COMJqkKYmlYM0iV6IuK/mbPyoLXJkPfT3bfcyZwPVA4trArFsWEE1Jb4XK8QhLflDMNen9
Gtd93THPX1C8RnkoOThQYq4TnLn9MAtgUOwOSyfCS5pnz/wqNfdsn+PP6ZpmRMnd5iRfTrudEWTR
tcn4D67GJNBSLiTq1F+POKZncnsJYXbqGHBRFLRXLjOoAf5YFsPFov8BHfcp6I/Q6CYqwAOYH68G
UBuXiwT5nPsB0maNL8o2SUOngVl4m5FcAK0yPnApXznTnvl3zLnV361qADEmEwztEogzjSafcc1E
G/VQT9eFrk23tSNCozWY6NW3nndYn/h+Ca2u5ljjQkM+mEIvaIVXlzpfmLN0cSWz6T5Dhp4vBsBc
ZYQWZF6hxc3kqHBphm7lqVv1cVdvE8zxrJAG/RUtbMbOFv56xfH0GaFWK9DjIlTOsRcct7drPGJF
23rkZmlPRhr+E51RbHm+PryIqlAcblNqV6H2Q2svXyJYVMScUgRWOQ+6J4IdbemnB/+3QxmDDyhs
xkVkoUYgB2izUOgao1zgdGcI24sY1vNvAyfn/d18TQ0/iuFR7PLUC+/AD0/ICJ5d1c8eYoVleXtG
6zbJzDKqgg1Q1AxfnHHrVYRASi0ipvNcoG4jhs+zXFVaTWVKVPn8YdVi96qcjMFo3j3MTJXjMPts
BnrI6YFfi61H3Yd2hHeDuO3py0OoT1vSPo8FiZ1uhEXmLPvZ6vn9jyJgX8QInHH4FiJt6a8lNNsh
wbJmcrQVtiUw2fiyes9+l8D/Fvlx1p1QeqXcoW9IO6ibsCrbkIQPkvsgqfRgKU0aud9vY/zIEqlx
1TjFP+iOABF3C0/SamOeYJufGm2Rgy6iVcATRqLJwErr439z1nigVEQ9bYJyswDZJqnecvNnteyN
XzZnv8LWdkbQUN8fPDB/lG5/UuPyH9AT4eyQaWJe85cuIEwm2JS78KlM7uy2Pb7LBdI15pNARTUB
/GchoXJyOeiXPa5rb2Erc2Qn+tmPGd17CPN3aTFq5TkA9o7e3cOxImJt4IkOBRRf9VHUYUAGbOdI
+U1dxDrpqnLLlEuQTSXoaRD/mE1Xn8sDE7emo5HN5XKgIfF1V+Gw7NRTX/yH/6dleLaFUzu+WgnM
Q4bCa+ODai/QuWXkSPFvliLBU+ecKoNPd9U8eUhI5qoCYTj1nLlMTl3fB2WWOx0yFnN8NG3ErF2i
ieBYS2SluUtdV459JPnXK5HdPr4llm6t6j5cQIpIVLDjjgpnc21hxEIMVqbxn0d9/EtF0v1FkJat
/2rBqi5SIj9/1MrIZuA9bYZ250YIG+yBDjUEMRCyhCYnl/CkGf1K/iXR2K6lB4Vmo5B/kNLoVBTu
3mivvvn123Y/LAd19asm5tRmaPy5RclyAfP6bFye3xXYC6OqZ75rTknIgGUprrhzi7v8dkxmG7Cq
8i/Y7KzJ87NE2GO5LsR5Tt59CbgoFp87/diQIcDBW+KIzhjQFkG2EBjS9NIBSPApXhaI28hgKUG/
VL7NQQYx8pKIskTlBdVzbHFNnzql8GntnaUfZwFe2rtf1LbIYaZTzghFlJuKbmFQAuc8kftp3/S1
wQNJz/WUWEOG+pyY4Qjc9XFexJw0ym8E7oxzkN79pyIITQSlWRJWzLz3X3nP0ds9BMH70dDjcGWX
ipw/OEGIeTqvyS5A47Mob/IirlXTiSd5tjsIOBLylpzXk0To8TGVJZo5kCj93v9777hIUgrhpTTE
q8+y3wfumKT62KKZHilxoFeVpPWhdOa4Vob58kpFeiaMYrnrhDfw4yScPf2OGkZU/a2us2uQpv22
ebMfPV0LaVc/JMq+hKIksyFMu3F69aaXeW0a/3wSRL4I73nzDAAngUUfvLOIBGo3DaQvsVb6V+Ka
qlIpzfD5UADq7j9Cw+kS5nV/6yqaFqcjpHnKYbrugwtE+qtIfqIaGoydFNnlhQpBBn3qd+XbVv62
5azzBj6On62EjJOM54WU1bH9mS4kvr/TNMvfAmXSD0IiOjELCUoqOo1JsFmuWRQu8AaU2o91x3Bf
6s2EQVk2XIRt3OO8pF6q5BTTWBW87nQ67ugkJ3LCtXI6owgLg+Jna/SOt2xoNmEzUW0kQ5H87vao
8wid3l8Se1IOlCcJf2po8qhTWF4MzhzSU7lkR/k/UNBmV/Dl1739PuyT0NK/B2O0w5W999fOVonr
S6KjaOoP9BLsSwmmx3ORIuTphXAf9Ajif/YFymXBcW6HAEqBNshDQBZK9w2lwX4beyRjomfGqUWP
tOqHrE+QjgcG1qsubthFx9ECzItIP4n1Y7mPSbUuKIeEl8tlb5im1fvR6eH0vvJOMtbaMCOgYI2N
ozMWEcEvVxAXNa3GlgKXPcT/q4LFSHzdx/jJi7LW9V5r1jQvd2qKGMcZ6D7wAqIGAWb0uyp/hqkr
pgl3qNcK2bn8XGx9zGNsX+PI+CW78KgX2wsUpJ3NIBU7aXX5EPf9FgPYdC0Ss5/ZE61fVFu2j/NH
QSs6EgdUAw1JHax7PJtlxyuDjVZ2JcSQtSUn71XLW6PyV39zRvlc4C3dO8MGI5YovaKkOWaH9VVE
WbtjIBLuBNGeOvCTxIf++k6gGOitZz6LftCJ/Kuw0XkixchoHmtwCNBgyUNH/21H+CVqVgDhqFIN
o13kKQj31fCLJHmVK3nacUdbjB4ZUjk8GTAuSRVHxQmPyZPCQEIA+YuA1Vhu8jNx7JTwX3/wokWg
IStbgurUVJ7Q8K8szgrSJNkpxCYWd5YWYJElvOz3JzV9rlaI40ixobid6QYjpODKOt1UOCrojYUk
qRjqrpNzvyEN7qQqqNecfNLY6JTJMNs8nUBfDM5Zjfw5gqbGNpEyGAQfsUBM+kzlfiZLU3+aIEJ4
3hardiZ4jleEjVyia9uuwfOE2YqyRyeIcqdhlJL50CbHe0j3Ugf8OkWLio7iXtmXN93wuV/7r+E2
YSq+9VVfaVmVpGei7FukwgpXFtOz/Sxc6j6oO6vHIU8DUo9vThqopvcAX58eBMwnv1InbSKW9T54
D3seNuFobwQr3Hf1NjnLg0HD7yLcFsz5TBgKWIkfZMUoQ7am97U/W24h2iglDx/fx/bGlDKnJOQ7
NzVctedLS7IuugpkznDm/+Hu89kZ9LBKlQcNi4hPXVxT8hMF7DzME7L6f2XgXdDlsSYRZqg9oI0q
+fE0BR6bVOednh91Wv8f9jyCqDUvS2hk3vPYaoq/9myKoNYSF9nRV8AA8Gvei9Bque/K6HLTZFIp
d6HnLqcxMCbc3rgslN8MaqpK/8n2KP1pJ37ozYZk3mFr7ii7yaBwCRKhBL1q51Ys6/2IB08154oy
zs8zN7AdQyp9ruETRJGIMn2POqx1simQoXNywIZXxBUlWkAoJXIZ1YrMmYMajJ09/0uAgzYB9OEX
wi3AlayQNWbbXBzjADA4sCPGG/wqEsVU2LCkOFuYA87hOxyOpN1wYCJzJKbYXSvLWl8CpT0A1YGm
gnyvsyxCFXcO0t/Lmohro9DdbjG4An0sK4L0pvSi573A1XhTccyOO1lgRMbUMZUEFQUaOzA9E7Eu
dVP57ezjtNKQfJEqJ18IZ3bvi1Bb59t/aECD7rlwodQs6t7rkRNF6UUrf0Be6qHkk9xumyQC/QnF
z09YSU7Jqr4Cy6qAuciq5xtW1HCm0hXHAL8ckCoBB/7wi+RGaJytFcuJkMVe/Sv/Acw9yvHrNoMA
3frfswBR3Kr57TYMv7oPWDb2nhfU9KsxOZH8QAlIpBFfe+JJIoOZgvwAExR61ax6QeLM7gi8VRSu
sbkfSufy4A3hEMueW/LRJ6jTB1BKsiNm2f/XGarUjhYcgWNIXiU9OKF78TdYyoLZ6jLGJpvXQPw=
`protect end_protected
