-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
a9SCVkKhIAtADq2yugJH5nGJYr4SIBjOj6XngDhTp/BkY15mAjt95gld8O2m84LBAE59PEIT+BmH
umItkIY91/nVSK1x14akDKZVuXvCYHWc+ShGyxeDORKJEkjD3fDR0ayaAiWHE9UxUdnDYvYnSw38
6E7tg96USWtJr8wURTPyeKTSsYA9OaLmr7wy2GGOCVcCJdddlpRqVaGRjnTOhuQLwS+OfURskYFr
Dyn/lmA9xKkLc1kbsYvnO3YtFtiesjiqWuhp9iTFydfjk9HMDaTxNFi9mciyl4y0/r8DiREyWGLZ
SG76nD/6K0pdaj/PbhRLbIYtCW8raDzMeb48kw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7024)
`protect data_block
jIoe18yfs0QflyKhTAxKHwDkc3TUBgMmcyDsmMeOlzNcXxCgiU6ZJ+94Vzg4RM9MhDH4t3fsErm1
USI94bm4u8ZeeOX6JNdiBkjHSMtMLWh6+cM6wXA1aA1k1mAIyL+hDZniHCtFRAmfCbrJsg+6Cr58
oTyspcAD6KoOlP9+mhpR4OE74SQw87HJmDk35DTzvdCaGj4yaFzsC4+HazKR+ZIKrGoc8BGTA/+q
q5zYsF/C8ywKSGV/cjbRZWO5aO7Ja1n2oLLwlRDbS7l6aqMA2VCfZu+2437bjjDtZqQLyqdM7NfO
SS8T8d+CAkPSiNscqpsP1xa+2xNzQGSaiBAYWluKSxmnrKDDsoRcez51ghQSLoJcH/Dlq2GZNLrU
F7qGYdCnP6pxdoRoUOxNs60B8yWo8haeTXz6GYh88RCS8KUHWHcNeMueKzo4JhjVpoGJjPsw7oAr
EW1zqHGH3Wv4j8HdM2brVzJ2YQE5ZtZb7aGIRc0060pLfcaDbquRUkYANARWAxQBO0xdPlG21xEe
w4xGE+yobCKusgOFa039E6fqxRrxS65BvM8NIBuZY+qNz9ATnxwsD781BAE33uj6O7C8lv3IYVer
mXVNivN0yvuvpzgCsK29ECD+skjBaZrvQvRZtaBQaKe0dYIYWHnSYcSa+f47po+uab4QWtIMbrXt
rfjKdIQ/wY3v0JSY+4ds4qmxMNRyrCP1MnuWgq20UJgZlY98oYYNiM3MA786WiAc7g+O/BIEYSGm
iG2xRhyu1ltL8/NSatR7/PTSuXPMzTA03oR46J3oZMFnc6O0F9LfjBtYBGFi3U3pb2X6QQJAnNFt
kR1arYhOontzdZN73xJjNGs76D6BcBMsYvhAQrVKSonyt5VMjtZhh4pMI1hk9aj02y9UWRh7nSHU
Lt7HVB6IZJ6hYJGX79+05diks6XM/Ehf8LAFM6mzUteH4CUS9o1P2QkycTlJlAG0bp9FI4lQh3Ya
op9MoCuyawJVabZAqGwKB9l743X2UCMOhu10nr7EHfULFJ/0VxeQqEutMqYtbo6w92tfOVYdpM5K
MyRV7BzTqCyjzlnhneGSYo1vaQW43rCa8/cNIulkejjd+UFElkoF/PrGR3QsRtTOpvaQ94x64vWE
TLcGZtUac0/mJm+jqzeG+5MyO3pTBvorVKYq5n4m2f9IZVHlwNm774qOF/LHFsarZwgIvs3tdzJA
4FKaioRcnfWYbPcP/GmHcazhT8CnT1IVuAkRH2Mk9LkLpY9H1X+VVsEvzqiqz7LSAx3wA/Cm2nvC
qkTZ6kb333l67C2S68wRBl/uirrUxuR1SqokIdFK2JVLAvIbmubUT50vQ65SbX/BEFAbkBAmCO/s
XtWAmpf44qWffPxo0QtaDWfv0JWk/zUK43uYDFAoKvg/WnIEqe2N70GKPl8L4FI/un7qxXFJhQ2f
OAHatZrOpOGy5yxQjJqDtGrvoF8280sjmodzS+1rgUJru2wKEl5OdT6Wt+Zl4qX8PGct7LldiL4E
g6qBOMjQMc4u4XleiQdCaObNVHjFvXYmCd4Jpr2IhM9UmtOm+Z2F0OE1c1P0/gYPloaqQ6FgMa5a
OY2uiEZnPyRiHJluhLRA9pUPuzsPAYMC84lTAaLEv2UzhLMhjXXbTuSanj8DtbuX/B7JXqokfj60
ibZ+RZKpYxhCQwBB6FPM/VJt6IAUv4HNupkAkNSfXhwim/Ly+ukZ83GTtSmfyITnzbNaoZdtPbTj
XmcXPi0p8masYR5/CrAjXAhjcHrJyIjtoFxSrhsoBq/w25l2QDguxpAM/kAa/KHkRfr2kGw+s+FE
WsZzPY321ruZoE5BGIVI8kHGJ6JmwRHiiCJ3BCToszeR9gXJ+Yh6Vf0gcnCMf2vBI5HAwj4z3lw/
pZuSQsY4laCoVu3rUQF+Nr1ULjR+xfBDeQoJQGBEtKaKwFjg+0lLlgrX2HBNXN92DkMSAkOxXF7N
6krkzi6NP5Cq3M5n7QaFrAuYPj8+DOJkN0ej70oppudhfwAeX5jykBmuzwp+I7mfpaUiVg4ITl0/
QzT00X++h1ZwMLYyh/dt5zKT7sDT0Vip5K2GdM1s5Xt8q1eBr+S4ny3fEENQwGmF3CSbI79PHG5e
b0smwN7+us1k0Vziq56KGG8QUp2O7VsrIPJONGS/ZPa4caNF37KTKOe/v/XylEMZZrQcdb1jgFFe
VxPlpGv7VaQALXlICPYw8vrZW6xCzNTchNSPNpOAnP7p4Gb2zQiWnBEesByM43JwipfnRgEeKZzC
ZRHwMPk06hLNnkLIa+XoehZyZpmHOtyzkb2Y1x7HC5R5IlPQgecPAIUXqCkRZ1SxyuJRdj0e0MTv
ywBW6SWa9H3FSmStz6jYp3efHAvBpXcyZ+tMxE6nTljTDxbILATtPkBByjoasxoYigh1VmrDdgXY
/sr5FN1iMsK4zbf7v2D1v8JyBwwsE/vcnVbxzVLtTyxckH2h1q11k8Yh3KuVGHH+esZDXZ6nQBU0
KzbqDmUic1hqQfNmNPuu/yeVxdfHM5Iq2yZY4bYLcgJ0M1FWwhHF9btu1Nl73vwkfNxpF+n9j6sR
bSDyGu7Kmexz3I5pYvUALk0t7+Ge4g5yhT8JxpTMuNQN99H0L1yJx2oP+qrZFJlCbgz3ih+FN0wR
/ieM+xLErRyQ1OzCdHHlwuxrOJqMJBn++pEDXij9jF6YLPMbAqLgY4D9nuHJuhKPGV1wHefSQ4Vk
ekTI+wWIG3hRbs4DXkHxAjbhtejv8D7QCFWqy+bujjEIJhaMp49GBzELpEiewC7jVG2cn0t0GEgX
EN7I7g11qYImzEdPHYrus5V/0gK9pmtSiGNA4wrlLvi3V6eWJRmF/7Bmmw9DvMOfCC/R1ZZbWscl
yhkwnVGGOnCJYqtj+7sIn0XOjWIB6w1KDtiCA8im2Bwyr9oNogGeSIyKXhb84EiKqB3vRBAvchRU
C/osE6YmBniIey8bFHeqLXTqfRVEJHT8xuoVQxRTvnVQqGrpoOPHEx67DIVW9+J3s6KS6rkXeILp
UT/6spBpM0UFJ0fEStWdkCC/Pvx6HBhH7FzwenelaBTuJqFMfEkiv38RXl3CGCkCgD4FSOXo4qJU
q/We9IMT41HITlJ+wP4My2he1bxcLTRYrge9O9+HuWzr3IQP7vKDKTDYyZwAFNtYWSvwBJQb7sFi
3E7qOGnnK+gFfLVr+Q0fgdy1atz9luVaLFXaaGBJMGZG51g26OsUwstvGRuLh37xox+gsvIOZR46
6DvGN3rN0SEvQiox/wVlt9xcY478Wf+7W8BtgIxXfT62pFsHtoxIDshUfM4R1l0MyKYwnV5mFi+u
HBbCNlCrRY8uuY8QSJ6trnfGbHbF5jnoukGWYi6eA+FyeP6Og68eWahiHWcDCoaPK0837OR88H9e
h36KdZC0jZghmTAfDaMbUhR+5ncqE6TUDirzDKVKhb0E8dKF8fV368o4ihdo/SNZrfIsPRTx2UDS
dAQ604Kjm7L+CAtNEIJZ/aUBvGApqhUzySCr0d3WwesEKhH3mGow3911RFALJA12+XB4YW/V758r
BtP81RHMkDb8vxzigHGtBDjgR8CMtrEXDsB3UEM35NuY0axFEGvnaoEMqctVK8278G6WsatTWmDG
5YrhGSZ7u0LmeFy3KM4BIa36TF2NaypNmIq/T0AG4B1YosS244C/6sx0U8jJLB/GOD1tewbjk60a
vAbg/2nzq54vWHu1TB7XVmLdZwhL8M7k5oNh96ISnB1tRfVAncgQPM+gyq65Z75/CyQHK2IxjYp/
Z5leMHXm7KueYdrFy3g6nr06tV6h7J049/kdk6UnUR0G316aKOt+L7wXJY5fYFjCV8k17lVcVIkA
BxMiBI5HUZAOuFwOYx13eKWPQLk5xlMTDHED9GpLhPtuTWlppcjrq6A8jTo6lsph0RNsCv8tqT3q
c6QDnDGuCh+OuzEl6+P3a85Hvx89UtxlT4COkWAAwJQfg2lzQm4zjHBxYa6h0XGgNrW0Ax23/3Cc
4qFF4M1o2o6dFe+ZEluxz2ia856yjay41onFIGg9izc0RuLdL22t1zP43zAqdpLbnk4cECbeHRkb
YWQclPUSSfylW8nZyRVUg/rjIhWeMV1PJITU63y4febFbYj+FojVQpt9hYwBP+v50SOeP9KLkNck
FeYVCPQR2sFLpTKcIDl8u5h4SafdSDVGFKi/+ZhjTfVkr5gZfG3vxjwy4ciOQInPb0u470f2p3xw
SBZRrrqgp8mDMj8023OGFjjbDth4/mHubKxjfd8iVahbNSEGToOJ6u6O28f/SiXKWya0QApIQM6V
aqNQPOKmLbM2kvTsn9SI1RYlV6WpXTEdx1hxvBb5AZLxB1h7xAzfOvK9cI+fuHftUeN0RZWdjBhc
+6+IIr3bvvrw+X+dD9yjWDMXIq4kGsrPC4LSjXqiGCZkTEn4MrQjPqiZjlSa8R1nPMrp2f/TIzIZ
GVsjD+2US+Z/v11Sg6REbF/BN4MiJkv8x3s/IoW3EHBD+GXkjSf6YV9QO8zWn75FR677Dw7786zt
rPWBLIxW7Cc7Kuy6HRrURCLaVlXTsg0Ee+qzgg+WIlsD/tFmld6+z1LW4Hbfnz17AEg0nOpNNQyE
mG23Oab153B45e+Eit74G4mPlpQ44G4bx2g218lt3CykBM6iQSQXTwYTIL4eVgkuXupPXTiRffy9
q9gousms1Reb1+Hg/9OfpZcNucTmDL9/KRZC/XKobsuXLKJFbaLeZrs5RtQA17vtAdzo04Jxjy8f
5J3ho3lo2Az7Aip+r7v1TxbXSaijWiFLRHwEAI9NWbo7rRm0LdDhs+KRPa0bRifTa8viMQcxmwmm
IvBm+BglS0RVW1RaLhMYxV3CTZnkLPn8e8Qzx+HxV3jOvSKABrkAj4WfWq7HWvFYZFo7RZF9O9Gn
HpJ5sr3pX8mtSXvJn9VSp8Z5h7GWNhs9OY+SFrkmZFiaLAC/RcvfS5+FLfs5biCwHIMdgPOXnOan
PX6RhIbvp5Ygf9qTEBS9uK75bev+ekgpUlYxOOS5XAIpPLtEsLqnrqLmDvkAEntCtVLnggJX8uTP
UrIsFnqr7qgronpG6xzxZ/KRxP2CNCf20AH7p+3Cx+eXkyNXZ/gytclfwXjKBD5oQ5Qn38L87MYT
rPKP815Ym1UfOMixX650fcf5SiRZJhykJwXj/Urxjpa/hdu6oGQpKZuTlt53TO21lArJN8zGJe2W
EOmPK7BPIPc/QiHrVLtlywy8vYAVb36TlhBkpHqLvexZKDdci2075Ym713nhLm4RDFSbN9nzKMCi
ZKzchqgNMuLna4ka/UdgEj37MM8g6mGaJfuRrXjlHG5yaXBsBGPBU76SoLnn92lnoVFFtRKTDSFc
z3w4DUn5tDWboALdWVNl+dLI18tJ0tYQ47jcslC3CcKC36XgsDH+t7OPvdKA7BPkxvt/y1oqGUBF
YsT8inU80/lShhsrcb90zPKNZsHHFfq7P5cGbAh1HUZLwk267bhokJ9FdKck1srvpg6INIQvs9NL
vann2pk6xo0s2x8R1DcZQkzVASxThLjrQboGbasgFScF3t5yP102M837rLm/fetE0HKHnjOLSYUG
vOdTP3e1QsGsd782Ohmc4OkSeOkH2O5PjURyilhcOD+Tjw7Wg2+Cx1RfcS5BeW8Ggj/wkXmwodUU
Mrfw2BCV/w/ArLful8pv2iQA0xXG+EDoE4RnqqHHOWqJMwbO1wz4x0DDIfjwkWYjNmqD7KSnhmCm
wbXwBPWMVW1/pSSflE6zL7B8+IWqb9SoffW4IYVCwGwiFJI3s+1Ku54I4FJOSfog/UiWgH72X79T
K9OcPONjo02BcCju2ak0aDIYh4GRPnzqjb4NVdPX8QGzhMRb4t/btrjx6ubJoKaw/slUmqedmlte
ThgsiPoPJsgPdGkFclCdTlLQXCcHF5NQ8nmx35rBZ33OOt7WAC/GQiTQpGPTModo4Xrh/vDtevl9
D2R2E+0oHB2r9ACNQm2vkSJ3Ug7upDD3aZ4yI7bR6lkpp2jzGfRlILtQEzu312iGnWCtP3uVep3f
OsL5OHMuCLPOiSoMTM6a3snXKB0nmoHsUHjz2EqAC169FgughgHBBT8+FfhW/QvYxAkk+BYFm3H1
5cxuS+Z1jMnUvXH+d9gL/kvwkTA7aGfvVKcCxeyUM9Ovrtn6picmeAAca1/AP8TnE3XbkR+LcIMj
TaPrUdURAfCOJ27ZRyH37y6TkJwOK4+tZWAD99/9WtBR8W8jnAUxO9IfFmM5QeitPf8JciKVbHA0
qLmf/BNZM6UDxv+AjvrEXSN2CtQ5TnCbyiNQ4UUt4ajfkFNeCsenIJ3LOHxJKmsWRykiZTwpBJ1l
vk3uwKW+PlPcDkgRXvDmIOYDFGNmVdRfXbr7nLzBQdAyze5Msgl/ydIl5pdV1rv9RyLwUJOH0ouh
deistJQdV7U/o8WFq8qveLqe7eGjjwlM1POyBc2nwffgxy2fMqUzvOlTrDfoB2FRrYvO/AxiayEa
s6K7bK7lKXQlqzuiZ6+HS0Ktu2SfM2k3/Q+W3NYOaXimvWcPwkg4ztaFNm2BSEK2DmeEH8I+dB/x
qyfUqEEdLOmZBcG6NpMK/d5EWzwILr7lFd665GnWyvTo83liXSMmsGMWdJMwF/y+RYjP4nvLlhdI
MszxvlY5vGLIbTeBHo3/8C1vjSuenxsh+ovBSs9XuRNlu3TC/vo0YLTgyhrNemNFCYUZ/3QHxiez
/iIgU9PyYH8WNLYwQkjbQ/+W7J4s4ZIhS1RCvK99Cp63MjE+9LpPRSa+T5nbQRWZ3dH8BNsRLiVO
Ce2g55X4lYV2vo1XVoUjyqEYNX016H2sOhNIKurK0bxyioal7jpli6vMCMs6gymeuTFLL3xD2sXV
YwUdtZ+UoHuUVEFE622sHbm/PcEQJaEAsynqop7gPidYkiBP41ZVy3oJa8DjJk7kIGJTfqyPHMzg
ZnxJzsXnyQFhO6/vbJ4sroYI+xT+UI/mIJx74ue9b9PWG/DCohWxakGTqn1M/o5Eze9mSioYdvsr
uR4dvIL35LNJDFLeW6A5/Z2Wt7Qn+fhEnCwR9CbV2MYHtG93DL4U214sj5MG4vaFFsyDojH0d9no
Rhqd3ieRsh/gG8DkNm5RIEok53p82GWD8XkIRKQ9vSp7kxLcjK/FiAZk1ucxORYprhSc9ht+eYah
ZSt/d0eH/X40+HShK05S6e3hzn4+rx4WKp/VX3pkrNr0qrLPIz81564XMS5ygtjKC3SRlHdbO95V
mfCuvwv7YTdmpvwQnotub0N/RBDIHaqKLvvI4u24kRzXmqti2/rgbIZgXYNSZsAur806mYv/6mnR
qPMofiUzvP7GevnXQkt5SSnaIzUpbqciLu5Id1KZNvQScPZgaIrtCJZGi0fJC7zhVjwyJOrZezsd
XEElWgPOwEuYzjIKeOtpojBJ0xY11R65e7ukY09HEiONQN+kMHl9X3CtwRUglcyqgtHEHbFDMOqO
y8kzSvd8GhmMYj4QUd1++H7LdYuo7bL1CDTZ3XecIi3Ar2NzcLtpTZLSeMcHbJRf6nHnpM3jClV+
8yeXVFJQM2BnaPIgWGP5/55Hg4Z+b0SOahMjo810dJArp9yER88h/iWZR4ZBZuHgEq9S8W2/l2oV
Rxmn6b7akWyovHIbQ79PAzYkdrbJ6ZD74avhOueUYb2FG17EtvVsHd2hC3M04pmaCc0l1Q7Ni8ST
XHmLhbru9wpuQ865Nf6LW8msKKgjHI1mlcJumAMAUbyy6BXqH87ufk2rEY8Erj7YrEVV0UuYmPHg
AqPTZPw2JSdrwXKyPLcE4Kopyq93QKMdkCC54ALuiCv3syQdjVBwoIDZDHDskUOOKJEY70dSqlCo
mKdKmwWlBnsXmuSOJJrmCCPSHYUm+Tov7floaHkdu4cXUnexJQLls6ffkreTGE+GQTJPlHUPK23C
8FHmZUnxtjArOMaXwAAeFeKT5ojzIfOr/4XuOggCkhzds40v+VRM9sk6Db33XrSlYBCU7GE+3Z5g
OcIQRyXKR9N3u9zRQKj1uGMqdBymB6/qFaTYuG45znUggBIHw3YYW2OKtYpgHg8WXzgYj/MPnTVv
pF6hyquC6pFUzq8M5hr9Ksh9jTeSIutmM18+HeGjFIq82Pltp+jk53tufG6r80SAxuel51fSJqFs
Q/dplUwKRxj5ePk/tu38rcQsY0FLkUV35JjZ05dES/Psv66cHh5tCokRIKYJYG6k3aaqAGJWsP6V
C4TQu9IYQD60EXI+AevW/cYDUpzD9uET5ZsJY+d6X061Fb/eKXI0pBbpFfl+AyIll+BPbqiPFUwx
WHKqEgDrVkQI1yHua4cOoEB77KEBXCHA4/Rzhhc9QY0FfIgSxG4H6LPUsIqDrPPh/Z1EvJDjLQrY
fFSKV0N2jqqb4blCDxqimo0hMgmDh8U+y5vwhdDH0D1IXOdGQ5qQa/9EFJpWsMhwaJqJtm/Sx2hL
9qSP7YRdEFW6aMLQTs/PzBV9G+hkLdxem43quu+VHd02X/8ifqBdMLaGM8Tzb5Nl5GpBrIATmRee
9KS3p2vl1OeFnckSQtqKmbCL4KyWQsgxKaZN5YGHVTs3KJgqmE0cnLGf0TbHQHw1ahZfQRfWhM77
dxh3/bK2zZ3HkumeUqlRSSVzXuuwpzy2hCPiEr++VYdZbviDczksze46LXX/mNZ0Du00VDPESONk
vMgtDsF1ibcLmj/k4vSShncFjUp/lZDXUFS9edxPA8pXxa+9o4XeuGzRBfWXfk19WWL0UsPceiYc
DNVV8Y2GiYhiF+faLntzOJVTIQknEucze6kT5msQ47EpWaKVHMlEqr9B2GNAcfgytbIStxR0bwl1
slofqM1ebYCcmBcTPWKGAxzyVS+mZRFHgtBwUkcs7F7dqMmjrqjCAnQz+oyxdMlxGp7BiEhjetdF
l5AQsuFhF/RjrhvZkjvd5gmTgSiOq5sa+HcA1fRss/aHhmA8X0N1Nd1ryUqLYREqQRPf+FqIj+un
TXTIxxRUol9qagH16cBVnN82i6cYIM8RO3WYS8yUuRMF83m/PEsjHUOtDV9vzPKtDiLQ0kgh+daa
hUJXLWHKp0eeIziYpfufmzMuQdvM/DwtLGkQsS/OQwS5wAyCS7HaqIM87VnUAffW05C7a3qnOMCy
WXOJ9IGJEuDKujaSwoLftZ8ffpxULkbUtOz1d7grD6Yx8jTtIJ6csDbcaqDWK8mdMxPIo7Bn5uAm
E8SHMOJiOepDQDnZctp7tq6fvuII/fnhOtsDdRMvuFO25PWN7cCgOSvCvNk5/QRvqcAooON7QBht
lL8CqUVZMO+QX1XNew==
`protect end_protected
