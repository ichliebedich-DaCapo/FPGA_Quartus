-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rlQp8oZNVWvWYrz88J7lG0I3S7cndJG4M1g67zo0KrCHPa7dwSgCmTO4mfXhm/PU8n8BB15yR8bJ
4093mcFJJoZm68xBhxIItuWKJyhr2tw94D2eLHSJBw0OetYCuww/b/0Tu7k4U5U7j01tWn2r/GdT
Tk/nLjmxFI705J9xsXgIUO2SIlN8gKOv3/TPN0EsZm07Bo2A2Asrbv/FrgnZ2XRfhGWjMRUbY/sX
W6/NJR5UE0tG96ZLA7+c9IRBFyT6RxxwJT1mz4ZlUSUksKPcTTEl19qmtq3njElEDAY2IQ8EsVVv
wNrPLoWbki60h8yNOWkum5rC7A1ulthtquFxNA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10144)
`protect data_block
gyb/bC6ZwBCKbtXRcF+kzHpFzf8g5xfrqujiSHxOpLcpesgaJXiCfaQ4CUWXv8nvPn1hw0pbP6oJ
osUZ8UYgbscJQmjX4K18zoBKs2qVqFzswLsa0RnquRGbElkTObSfLpjuJyNxM2mfg0WV54x+R280
9eyueQbYI7LONDvAlVCBcOIlYoldIE4vbA3U2D2/KTDsxLkpi6ppwqwNMxdtbAOSlPRGrIM28tqc
fh/ca/6rkBgt8JMf/9i7wOe7d6niuryWhgfLmPVJMKLaiIsCjcr8hkpEDWAZn+B2e8Y5FkEgAbWk
VuVFexEwHX9+S2FFVpExLuBzEFn04hFHZVFAWrtmtfDqslMvSUD8zgZe/ZPrgLb9dBPaqTRXzg3T
pm+w+zHAqE6aGL2LOdN+Sg0tCb/XkLqtlw2SHI27OhiLt4HMcBbWrSgVcWPjQt3OQyi1HI2lzPTk
8Y4yCfJsQ+IJcw8YqpQb4WqjtdOeEw8OU2plrCuLN+vmfL7FcfisoZHSfjv6R7SaW83tpqlTOCvz
lZYaM6U0JxjW4LcJbFHaVOxxkKe0VJ5L9U3Jzkm9bdkbdG9c3TtRkDNfEOrvrbBmcayI1tLspbdn
9yClDUs1tUsXWyMlLJYsQQJ62MNz6Qz9ECN6YBpgh+ABllniKqh9H//imCqE0qX3qN90EYjiyAoD
ne8fqEWdceprhf72xs8SfKeniKMuZbFHnocZEgJCER3Q/qtryI7t624LmVfDUDAgtFfZ0TZc90C5
q0T37wIkuSJdKTOMAcV/UZQLlyHdBj02xiwuZyBeu3DI3NO74TN23bACzt5CQDU2pGjh7PtLNRhC
CfKV7d8zdVh1hjx2AZDVd3XkJnYdLBFDULuq2lMMss3r/kyZUk4I6YNXW64+z/whj2+Tow4zZk8Z
wRgvl0YzP12bB2MbSB0JpvOaanXpB85hfXSCQWyBH7ieG8CyUjbVbT0JEhJl7upgAKf/ySwkmBS1
YNIMnPTZW+D5feJgEYIi/3HFwwBD+GoRWpWqrbYk978yDm8j8qvR4mMsmjkBLEvb7ls5ROes5L7s
T1cd+tODPm6WIrnO48kSPYo9Ban8d0sHYC6dJY+Ja242T5sjFMpVsCtA2WYXKKlRNpHMcSaw6cbX
DdVo/OxSaDx+8/DRhKvLDtlwXBYm7+aIcqaAuWyAmlvlAuT+bATs53fsQEsyQ9ySPFrleqYMl5cO
Csy4jKoT8IhdDC0bN2QJme2AQrkVSsqenl5Rr1CE4gihGF+DjtBU3eR7NjlCye0pductsYk7eYCV
7v7OSbZPzzfOsdkaaLPvk/ls74SF+I9YEfMTeg4a9m8ckWbRx9ZukA+AZ7m4ZmzAey8paT/x/Fix
AHioOmTdyIg6LO0qGjGcLzsDqapY5IS1WJ9t50cbJr0+JAG2rK0XLaYFVfQ077Tka/0Q022/hCMP
X0qpJV3Pvsqv2m6MmwBFu6zFbEgqP+13mLLJI/YzFAjfTUDdLdBFQaFK1UefcKi4wBu5wO4wMqd2
b6GnMSzRW/ngB68yQ9VNHuTFHj0R7Q/19SFTM7JfUTUfnCyckP7AOzqgmKQ0HQxZ7GTgCWhEeupP
bpLjkYzr9vK+dkxEyVgQ4EvOHasm70IZ7lGIOs9JHUD/08cSpMA2pc8tKgo340RNPT+0T8+H9Cbc
9tmcMP/IY5Ehk+xIpozdpqGWVdZILhFDJZbctrwXNE89vSzqw4x7JQVvnODn1cuVjcmgeif68yjY
Fsre6xiMiqvh7y1PW0ebr5ImCNpEiER3kjdFMFyzLKvRykc4+7m7yZWlueCO2QrusiH06+XnMAp0
qEG0I1QfdV4Mue0TgS45XfbgZud3BLvLo4NGnrFwlYaQQa8tmRpJkkod8AUxNdQebT5fNubH9V6+
P9TYBCNj4ArYBC3KFviVYCTLJNfvKbYc7ZPLynvAa4drfyJBluX2FD2Jyi7C5B647LllGLUFMMlz
Rt9BoI5ESb/ufpGA3PaQ+7uZS65wftNIeCmJYbsf1HJeiR9QsYS1vVYbNbJFvIaGRezBRr+d33Ql
hQUESje+ZRuvjK/hPIevFNgIdAK+j98zCur/2d4bn6+QJxlhLqbkC0e46+0+przqcII+xAJNlu4L
YSmV0rPayUc6DNRkXXWImIev6Ki57CyFStk2buVlFiIfLmbpa3cALtWiomKlX/Vav8RZwRm9uGdJ
KrAMRY6T/ZbeV8Rj345v5T+tjRWob4QHxgxTvZzf9ppx7q8Hu3hPvrR1GiFtIVwFrBhm1OnUdqS/
7tyE7vKZyha9IzxY8XOv9WwbHfWS1xcGKV+5WuE4/GYNijNX50Hnd5fdU/H8LIp4iyHtRYeux9dr
2tuJ7Dmg/hghcO13Zi1GvYTog3P5pQ3g+jRBFuOQ9yLetxi26/ywMumRNb0FfAKC9siht9G6g8lC
vA+ipcWHJsnGJQBfV1UI/wkQ6K8o7oXvy4WtBF+sGYjhmFlMJHupYEM/YCuM6gPsfNYu/Y5t+zv/
NB2hIJrPBIOMiO7HL37yWO8h2XZF8l47WuVqTGT6xF9Qp9+fN9eXYdGlux8d8L0qeFGSE1oK7Eb9
m3cm9zCaxRTm6JB6WNGDEpKzDVRnCMktq7HKK+y3bkGkjIYGL89nOPg9z9kY5MAqkyzvnG2RTO1Q
E7SbiZdVTTMPA9ttW+MYyVpbyOMsWLnXnvUQ9EslMljbUL8NvUnU9eDXOw3KW093m4XfY179c+mD
x1dyzb+091uNnK+cYSC3U48FVY4Eog0QIEB5ObVqRUIJ2ybKUV3M/5Tq4ztSNgjwywFQ5G/x9Cqq
TAWvTDlQ0ySVDKXDbdvpkmGgEmgskUGVBn9b3n4m7pINMJRPvhSAiTm69M4D1Ad/ptDDZZ4rI48M
QD4+AlJR9XKXf1fmnA29kvpPGEjmystaWzvWQMxbAvtw1u5T/cOZzD4FxCRogXv+UvdCt6Qpf74Q
GL0n//ojPf4tgQY28oXBedbRXVp5/kog+Owy0O9v+h8ZOFihp9aom0G5tJeDc60BQ/8PEKK6kggN
5KcmoA+6cJ88n9WJzPmvrVOf5NUZcqJtXqIZArEqUFTnCUST9v4uZ99/vPhAweOSP2wWZ5aLcKt8
KdMK58H1tUOP0f0XVZLtXO1MIY5tNpkJQjMpfhiz10HnJ8zwi5wvknRHTZ9mQc+2+Vi1WSrCSRcl
S9t6M5Q2PNxjBxifxQXKozNA9iRu+HOTE0NIfmqCo4tpiv6y/mZMytUh/KiJhMs2UcA+S2nuLv5O
3xxQcaQHtbhsMc8NaSXqfP8CpyGq98szPjbst9CLNhwQU/YOURsi9yUdYufjD/akfKMzLZjQtT1i
PUVvgzjxi6P0Fu1gNZDZ0RyV5aPpmtyZUnGnAFC5isUKgTOS+kiadouURdJxy8RWR7IybzNbeUb3
PcOr5/4ffZpzKKo0vgLsonrPbcI3QNLMBFOj+dDE883gClIMc69OlAxW0kBFUi37K4L2kLU4qkIv
slLbNLBqNd2c/GHxFRXFavVHuuf8D0Z4DFy1kc/13l1h+FUv8dBSTCAw57w0r6jTIVh96cv8oL5U
6m/wwq91uygsTPR1r7lD4rguhAcvspPDjR92eitJffEZCe16CAG82CNgzgyUK71BcqGWl30ZI0sA
Ebt0cUmg34iTzFBo85Kc2/3UYZUKVBEvcQPwu2xFPd5eIfWJz4LJ9B75mDZTxFpvGQugcV134+ms
oqtPrHS92v3/yHjWs1+bq93p1h1PKrgaHZcT90/M8SsM2q1hdJmf3rscS7G18FB/453WTtTSd/S8
0n8Tbi49wDXAW5Kd4zaPz7E1gs9TiKLih/lMgAEKeU8TD6A/G0pHy9RdmWxoomTobSWqCHc8cvYU
3csWJX3FzA58mXvL5r8m4CG6Y1io4TM1RfvO+lEjWt5nP9k0SKjl+W9MVu4UjyRMIIBptsAFZnuV
d0AFcAn1Hxz4PDTgC4VuAuolHWeXPRxAxKU/8uZhOhcYCxisR9541mU3L5Z2tMBuCUT95wL3+SL5
Pro5FX5ltnWBjsW8p7UfUgJ9JyABxf93ILEB9ImOgO0WAgmeAp3yd8r+FNY+62540cOOBOThZUbt
CIsn1zV8YqLIwXPkWgjKLfXYfcrSERuMB+XOy8jLCuUkgYgUipOlmkiYPVvQ2QAoNXZu/9OqxnvL
FJKRqRvyrVYWNtnqm5eE4aozdwGV/Ab6hMCWUUCWH1oDlZ74dlAAPDN+Ivc72/ka5pULYAslgzb/
gUxcx4FhtN225VsmXZziBoIYjhkKVtXlKXo1os7ZA27Dh50SXOH6TAhZ9Y2nfnObNuXEhzLlUK4U
50yUtbAaD7cxhYT2rnJ7eqJcshiXow6cWyX/NQyIiRVMwFbpnVBUkU3NsU8OotmU8NTYEWVYTY45
SIpKte7OdaLCZtihPFvLH7XajCEv8aI6kjASjfYRsWgG+OwJiMzBItsCjE1Iv8/jSedATnBnyrHD
RUSzrv9GzIwbDs6f8zzetSvuKNjkRr+zd8W0S9NqNmwLUv1Ylg6jVvHHxUzMJxdHHfjs+iEJX1oe
/0qcx20mc5jCtJX68EwwoeKj9g5wZ5g/0LHk9G5/891dw3xCwxfL3U+H9Kc5KuLoAPzCaTPWXICc
usPRa4gb+fRQDbojxJWcVUWhZpZpAk3jfP/WcgRmkdV8kCeFYgbM1n3tnd6oApVzrwuXTBiZMTPh
6G5JYv4qCF8UMuYWmYPGKIz+pcX5tGlmR77AfV4R8Knk7BUpHcY2kWkBdahJQXX5mYIZ212GjS/4
LLpfWLA0s+JAZa7Y4La+ZTSis9m/72XKBUbPharGF33Xxrv/6+MtUIFpYfmtqMCSbjI+XCt/HFlJ
hdJ0ZhcWdhp1XJm4pymk2QYXVtU48T/tkqRVT3gsqfbbCouoYRI12RJEmgDlM8iMeVD2GRzlpJYJ
PQDtkXnAFV3xUv9e4Y+Q452Lm7vTGxWDdLxge6OPzKzU+ISuufcvloEf8Ii1r0X8gIcHejkDLith
iV03zbLdoHgYsO7ckk09GB1cr2/ZvqpAHKoALJQ0IbZ588K536swplpWaxwmvW1Rb00IgqUURRbe
F8j3t86m8uTUQgwM4jHIZMAhl54wbBEIv+w+LXzl7pustEm23/Z9x6+9U927/Ob9v0O/49TXb6op
9qZl6x90tgSmpdEhJrtpMI0LWpJa8CzQVfLbhtrVDmAaod0tV/3mXjD0kvIHjWS0ABaduF/l2Pce
/aG6xp2gVOlFiXX31lFX/4S/s2Ofc3C+M3ASVX9k1r7V0mrSMShYUZELR5OTmhICcxhSxogGcZHv
S3xZtw0SqnMVVm+uOBrAfww0NDOXhn63RP0GxwdNxVWC1m+Eob2gF1m+xmiIBctYXMBqbLv9NI5s
7yMYVair218sVLQ1En6/HWympS+9UyZMF5wmitRsxWyxx6HRX6BzUoannmxEkFtJQI+TNYwboMog
hxxQ96Tox4RFnx4s0zZllvSxMO1l6Z5N85nh77ooEYelyhkfRRXtsBU38xVWALILQsUhv9jTii8V
dKG0QIgxEvdXAFvhKpH1XZa3hgtNcRFLFv671wGtEkiULfbveD257mYRPpzGgJHJNNFvxU6QGZQk
603Qi6tcM5dzLQG/0SKCNyni8y0AccOgzYqu4J9DKwYAJ07t5nRXJIdMkNqJb/RF2cnNgKik2nNY
VuHEdnTkNcHRJs6sdrb1xBOq4FKDWwovZNLXv6dkUBK7c7APvf2mwe0W1z8TZVXVOJul4uKeewBO
VsINt7NPW6ddwzBl0Dx/TR8Nu4X8fm9BSrIsozpj5oOcgEfwX8/9/gI018YtW77kXjq4wm/wmh8I
DMy4offqt6pMcsEVcsONkm+U5lSoLvQVxQXV6Oh3f6r3i0bWJWcMF08AgFTixmxZkteFR0J/yWyQ
iq6Y4ft95yAKttIwhe0gDhElPsf8GcnUJMA/g4G11amyhW4ADvJGA1tEuXqBSL5QVqH8PHjv/XfO
13G0aqOwOq2+EQZMFe+vzjzhULZsYyiCBvgFgAOEiqp1pKDCA03F9yteBcVUGZIKoLTq74VvpT7x
wcdx+jV0Z9ynUXN7gMjd2PE83pGS3FCVWkFe/1mQ8ON+/UX3oAMQrWJLWvhr156ufyWrp+VNGAS6
Ve+ZG1l4vKY6wezA5hB4aAPDFDWA0mBD5Ur4vxPwRhv8qwvwsRpWvLrpw/Q+K/HSM6O732cdXYSa
gifi3THnFp68QaDtBq2mL8dLDm1krXd3PKQq8n689D5krUyVCvG+fWIYE7myAKRZlN14BGIiOQe5
840v/y9kl3ZaKyASTyqLBlPx+HVEAP/SKILHxGW6f9oNpAMHeRxXQfVgAiiaMffqA8c17NRdnbur
RxBRri4z/cgKO0qsoPkzGdERPIyTYkvJKoaVTDjDMG2At9Ak7Dt8aS+rawWXSy7LF1I2hRrUkci4
HTxAvpvwYjqsZKrNJCWnt9TYLpsAFOmku2b4D358wHXcMMqY6RbItxi1YnYQpngkpeANObfTmdE/
uO7CiPFl7GoW22fHT/m4zunRlFvehVfYGMGE5Z5zfeISPRskeYWe5lf53Ru5zGLGCR7RxMiYw3mK
QN0ZU/FQJqt0gnSb5hsEM6mqoZN+myJbqA/5toTjayJfxBQllXgpmWxtox/u857HXTxdX4s8yY3n
EtFmA8pqsIWyKjNSSFIJf8c3jh55jx20pNteU98RQjrzbt33X//0dA0zVqSHtr0KfQoeVailo/3u
zlWP6hQFUqZUFazcEtnqyBINN9j/ECWCwdwQDjchWWTB5ucLCyEKixIMIFgas8W1VA/Clu12b3q+
Jt63ak7tPfpzlxCJSbXsHMXbQUHQtB533xm1AO3KzN598oZWGZvlv5G5HXObaO+CNeJAzrzE/VjO
xZ9/yn8TbFu2rX36JtUy9JGMH0XghRLW6rEcXRpjfuEX/OEvgsBuwpSsll5yU/SmXp1UmTS9M9Dd
x85qkXiy9Au/zUDZ6bTzpvcHH8gEDVUl8XJa+BLqKyVmruwW6Ay96er47j1o3BY1D1UmxJ7ZmgBM
5pLtXs6LFqXLZeU1GXknVev/kwIitZ3ot3N/ZGlUmuG5YvAH/b0YW++zkSUXCAXOnY4slE4nzn40
guIFh8PUWfJmtpWOICDAkUeoWoeB2FnBiNiS+dmkIOIQxPErEDYKEHlTtVU5KO6RlbBKhoyxsFXN
vs7g9fyi9L2B0Trl305RLcECUECzNuH2dAl60yKOmXaPZC6gualrDS+iq9mAZQVVkQM9zrrNLXLN
K/DWfrQQaK61ElH4s/V2PeEmqdiLrJE8XvPsrBeQD0ALF0TOcnMMqjfFrkPbfyku5wqzWmuqdikl
EXUVxlS8dh2VgrB0FA553TQYhz4SFJ7VaRv7z3IYRwCCaBx7DO9VF6OG8/0c1I8YSglSdQVmoveD
o2ZCOGcE24C7IiIaWG/ucw38TZEckfS8dFY9B6LsGklXXHAhNL0zIoIFdsoE34bf2SrqYXj3YbaP
7R0hY+a8YeRqk0j1FSMrkDn005JdUUrgwLrCw+qqET4rc7c+D9mzUb9rfs5YZAOLs1b9dvLadNCd
G5uECqxofFCaS/EP3aK0zRMn7y38Ll6Gqu5GCo13f6LnoflMoO4vSTiTTOEGoeRGukV5R/63H7tA
2yl0CTqJ1YE5ngBt+rZdxZs3SdE6koSlTxJ0DZSnIAWRVO55ze9DOht4koBV16O5KSEkL9XaXm06
CoLztDJX5nvpkyvk5drIWG7lbvZeh+JFzCmAFXkHDL9RZa24se9vi87TUqg8dEuEzL13oiqACcob
dSGKF6A9j5Wpb6p/i5oVROmoWTJpAOV45OG4LyUZ5WFsfqQPdkgsdsneDK6RVsMP1UCkr0qGKuP2
8bvdxp2S5/xwzX93CiKNBEq9J+rwavzlsgdSPYdG8qkSBunKG2hPcfnN09/SDu4F3msZwPaMi/kp
I7xRGD49mKdgB5M84I9IOrQqMzWR2wW6kebR6Mok1XghBn1UDQHusLRiTRZln4R0ijLjbozfrW7v
2k7u8siE4CTK4Ddk24yWFOYVj37QASNMYmKIagodGz6RQT5KeejWrKr7UlViwayJcFA5svShR897
W+bikuFuaaF8Zs89Pu+HW2eMmt7fbZdVlT3OqxQN2PvPrknmkfUQT1aVNScYHlY693Um8MpYNNYG
bx0TyfGA86Xxmx7S3D/SPXtwD5NrcPjr9wqXjB/WEyZ8MsiWkMwzLdl/XK4i8Um1GnNIR+hN8sLC
9uoj8r3a5pzGQfTHFLpTaITRIvvL5o1pmNlRdV5Qd5J5HBgYqO/+gfOuJkoukkFeiYZEtbhwHoi4
/Aikg5vl2hiHD+SiYo0XRCIx4W6rMPGNgU0qViYm6gWQoDHPy+/ILEckpD03575z4eTB7lNDcWIn
vnbUTjlXyM0B5/s5hW8E2HRfJnB9CaWWeRSteivmxJxyXO0RMwksHS8EVWs6VP9xXoT0Op+X197o
hEAhVb0w06AgMmgUDPrC9PpSzDV4N58K8GCKuoOBx/SAM7SJVB3SnpiOXYplE+OtgrCxcJDOL+I0
16y/HIe+caNWLdwEKNIV7pMmzJ/HoiHXp/LZV3AkNLTvkyQ4/OGUXTmU0QYn9zhT/rOaw8fquPz0
JphwyEh8tH6TmuI9mLybdgYx2OytNroGlnSENKB8UPGI6XO6lQV2qoXEQ4arMzd2cbTHV31tc7eD
8sLd1tpT9FmA+eHbcqXUKEY5P4wl2cr4l+nWnE93ByeyPe9jQdTXpivLmMMhtXSHMFtZbAvOqbmx
T6GyytOp5bLgQo9CmS753yTBYSWzhS7sRn2kpArC9HyBuFOyK1iodH12tVwi+zT+8HjFPYPKIBaj
Wv6+Pg6vaReIkMoSNcW+NjBfnm99Nj0F/Is3/3J1lXZ6k0FeTdrAGTpJgS4li2iWe1k3HNVfc/D1
pIS5Ke3rx+hjiXzwkfOfL33rTnfx84LbOIUE2u7MhPJzATDwJXdnIqELPpcngvoP13ruvVtf9xMg
YAkoian+5f76BV/zu1e7GomYSU9+p+MSSL52260qlCkYGaQ4iAMwa2C/Wkk8s6XN2l/LXuesncRz
2UTNlfbb9GtzEprHhwaHJeyV5XaGABztMb3+9nQqHCwoa2JYtZYjWWY4qR311itgFFSC0h3mRvKe
OOXu4QAQl7fyO7LsPBqB2gvAsmc7CL38a3L/sMVNh633c0Ei6tjg+GFZeiJMdXdps0rLuxR02ZA0
l0oil6uDT/Ao1TwWUn2XpGKPqHWz7sLOKSf21F+El28duIXfFctBM/SZHi9/x3lB0H/XlXb7gygP
NzvC1nFxVr8aodg0jOnu001MJizpknWoNXgPkTRoF3kqTiEivk215ipxd53XlTCIsDMYlCAadUXj
Q2QeOk0uYFrVTFlK+sg4K5NgEfPQNkobnNgDZBVIiTLDrkTUhzAxGX0e4juBEgGWwIm3RPai3gBf
tFfFUyHdABnMpRDjjhP/FimAcQmQE1WjZJq6RS37gHrayaFvJW5T67LL+SiCsGa0g2R83+SNuami
vnvrccLeFv1UzoHv1UgalUSD4ruDe6XtZiyXdaLIW40qF67yFwb/LzzzSD/RFXYQIqtDbHYsokY0
+rQT5JIYPlEWZsBg/aVp8xpctdOhrHrEtwOmYPvp2fBh7gcuNWqypc0IRKBEBnbVKss/ZULC8+mf
kcSWdwxhhRnHrp0DaIVpFZZqZFeGrJzuIUNe3iyRPT6wLsAOy8xAbnDuOKcBg3xmbv1/2k1IbSp3
YgAeriO6gqqPz/lY8eia7i763r7lxNKl5+glbWPZKA7SR7qYxl1cu1MI0nIrU4bDclnZ1AS2tRi6
f2hBE0wc2w8U+BZPEP7E0+qKw/IPDIyPuGov2taadBwMS5xVjIn/li452yjlXfqov3HkW0qS2c4x
6Yj9GVfTSO+oMIGGiN++ns4UBBWbziIJjBTSc4vSirbtL6sEtnGIKvGzABT3ZW7HjALvW0kADQmR
3W/+g6FeH2I8AShx/+tQUM9OLoc4YUMsMGNkSIhH9JbVVfQYU03TfTdx8A+kUz2sAYqsasrGQLEH
KKhkqmDDBt+KrGKFLH+FCqQuyqJXt2sS0A3lw06ewQR2HEFzX3bKhEarY+nsreefcUPPVumoOy99
XVMczmntA3VStMOuI4kkcmO+rk9su8pJr1LflzD+u+rbgGtYVsDCyxXenCuReTrKS62Y199bFaCb
54IcmwOa1cKsZ4E5Ksr09HZP0aBz64x68yuY4zYX6CHByBcSsIfKpIH/kEgzLYtNDP1Md1U/IJy4
5NdKx1pcOr1J2mZKq+SW/4NbiyEgac/Knyn2h+dq+nlKKUjDJv4n4mhhvlVEgGvS7HO3P4XLes/j
OqAKCy3LPEfuxhM0A4IhLLSqIBvW/m8jqIcluk+LhYP9Cwokr0dupgSOh3ZRXi6rl0HGzQa6RLyV
0UlhmNHLwmJVLihQeFOe7Mml7uogExjt1CSEDdvwFzRGHVpxaNLeG99oMxFgMWjKMW42NxzcS07e
FdlNegeEsI8rLYEICGfrn70rQdlOGfDmK8TW/He5O5Bsze+x1wmTqR47NGdFZyhE0e1ZezQ8B6xC
SLax2NFh+X1hwxOZQJwSkSg759jaXTgwwhusZylZNF7VGhOJHZEBaOgWUgNQEuviYKBgKomorcNT
jJNp2gAtxt6CWTCuIgwrSXc2cEcHiQpH7B+1xi231o5MvV6NGhlhkQZ7ATsssdY6umQ1YeWADtoc
2KWxOVOwRK4UjWZyxm7MD5HiYpFO9ONwyjWU/GbhIu5zAZ4gpVYaQD0ToG9ajvkd8ESwNVpqik2D
JXrPRO9dabQ4ksPq5JAZa//4bLvCg7wf5FKVkJfaK/SOFMMpffcAqZhicESo00n3xeS3LXCg8WQ4
XUT5iX5uwWWgwxeNnI71rimQJOfAEBI/zyh9clEY0ALqL+LD1hFSAv8MmkWTsuD83AtkSEqgY/d9
D1Eeav+5A+ohSwQPQz7gWbkU3j7NR3Llh/BSSmruVKoCn5snDW8GPENZAiYnOJgFN489nYwjtyk2
o3uyfcJaxiviMaidmoG2Dija6ySfXNWvhub0OtkbH1Ls39o0BRRt4Axc0A19j0NSqrjt3ouZpOhM
oFyzcAYs7z6y/bTxgmq0SAs4DSPSAUbI+R2JxwWONiRAzJavTZh96QL9nDfDZprm70BBlvTpO9xQ
AaTg1BhqCETOOGCxVOB13dk5WsJP8BsVuLQIruD6zaM5Y+7O5QT4h0VKJW+KjRQR6JZgpmIsqCkN
E3gBKyNdER2lSKDB8xezjeEhMcuSaeNyhG5SP65foCZ8lQH2Xa2DydM6RS/ZoiLhDfv1rrkaMzmn
LnP1X1MqlqrKYKeyj7gdQdXPhlVLfZjHuhGll0L7vwdcDx62MxRXSJHERsJROEyTgYbFHDQEsLD3
zP5kaPXUdh3WUuBH1eCN6tK+BROdGx8BwDbeuXroNyixn12jDF2xHrrTHh0eKMTkDWZiKDdNAGSN
uNidqc9VG4fKZmae5SGjw0y8LNejHEUTk5h0FRIb4alGIk49oy0G3qIyXu9Q+DE+l/GDgIcXRh+M
aBwsnFVOONzosIe++gyt5vbwftzuvO4bRtP5vAocSASqlQX7BQxddqGgjLFVShy6hyElwFuIlha+
CYkPVQDsmDZTIx7BBlr4S0BB2e7ljD+QnvOZa3IBSci/UijWGCQdK+eAA5aWEvYeIsSGlm+fdLjl
YxdjTbWOMwz2tuHvy5IPUd2fdzjBV6CNc7jeKNM8+j6Fr/8wxEEycSyo4Y7YZnGUTJzD6TTeMm4z
31MuJc6CYcAuJlcmFbEL8N1AW0lZtDUHRpfjj2qJDk/tDi+N0Pc2YJHjpmfFuMd07+dd6Eit3wgj
/zlFYpe/nNzRurEJKmoKd3UShUJsTUfRhRL5Mja/PyQsbvbt1eyy4BUf+yz/hyA65/bki8QUBv+1
j4cY88XaQMJge7ZXmlbtZ84JPaSlff+ojBEefg140lthgOcloasQaRBoFE+0hvVN+upToYp2IjRU
JNxE3nBi62h3nj9xjn5Yhn1CyB+Z1eSYWiKEwxEVQtPym9CycghR1DHESWPX5wJJ/6eUg7/Tg0VT
DlvJACMPlEUPBnCGKOEWsaBm0K51fRLMnQ7/joRljRqTuLXYeK7b6l3aHvQvy8Sig+N5SEBQfV1m
ewpDSbABVSD17hWAEIr468iLb4TFzrq64veF7uVlNehIPTw0evNQQsaXLiPuJ6JPjMPsixKlI3Zp
Y2h7wyIr1KIR+ry0/4Z/E53dIv067VseXb9pxN/gqxRnK2bTG7kggxZhf/zq6n1XY/1umgGnhaWP
+88uAdbzkl4UxOW4ff4E8oTLFEb/xb2WJ3egKfv3ns87Qtm46uFh/p5LpK8JcQY8VF1rG+7J25su
SMvoxMb0MYaY53IU7piTqDZ+6yCtACMDSvrKMT/iNTd3bab9fYQDxeKxVVyLIbgYodvqsTgxhuIp
sIrtpYuYnAeg4OEhHULEXDY9lpV/Tw9THONOHFKpTwgeUZW9zZ7s023dfUDhAM7za0ZHIkqKTmhE
9MJwKnezynWCS/f8zp+1LiEhteRbUQ7Fq+VKdg7njVe0WjJNYtuY46d+Hgul3dw9izqpQEu3dv9U
8/UsA4+N42ogr8F6+zxLDqOrksION8H++nI0zM38F+78PULY6SqwuwiiijkjiTgXG+9NaB4lc3dz
Js0D+SvwNb/E1jxNLKX7PGEk30PdkYS4CgRU/7b15rbd73oVcXLQjwsEVLZc7x6m4rhzvftK/3YM
6tP20NniXOhNxLa+ewwnPL+hESikUzGrBAKgSHlFwyIjVJBjLnybZk+L6IJTeCDnnqMVX9LxD9Rx
s+oUka3Yg0AQDrpfkEq9iXB0xrNM4lQtrvEX3Yjkz9uySjaGOYYBY0rxx0ebQsyNSTQHPwgf+I4v
n5Yi7eXdZoVtjzKOLwv3LIV+X369HBCBK2EI2NXRsmAy0GOPA+m5bXvo2uZmu7pALYERyHcBIjhT
zfNyDmfc9BzpUnoT3xfm6NJR8L3aYwVXgWiQlh/HHr6KXeV9xVnQNxj1C9TaM5l2jpvzV2ebNYLJ
ECTgVCsp9/QIeQ3grxXIZHJH6iYJTJyYmEJn+siwAU1LFSt6A5RxYd7mHim3TbCHwLyDf2hrOMnm
J0bxuFh2BDmkWbAB+q1SYBBG4enTeakY0FhzrzafT96a/ThBj5HRM5MiX8XS5tuCsKsteVGmGFIn
wN+3MZzUwlNnW+J4HFA6Df7y8tzVlH8c2Bxcfszjj8tMcmkY1Im5cxb7TvwZjNYDPnoNUEI+hZBg
bHiL4W6c5ehkobebwh5QGJsH7MEuxlmaMgockCXoPp5Eo+tvHUqPLjuX72N/u7pzH5kEQSZsA4Mt
6pdME4jy81NXaV16RyM1xbipAmp8uEelqYYfqQOGjHFzTn8ZCLBsTTnimtZ7GbxSgnQQkfavRA==
`protect end_protected
