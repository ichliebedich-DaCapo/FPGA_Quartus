-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OeBY4B3mFV9VZI6wWHxzFohesx/sGQ8TBYsXJemsp2XY2TBIw7wT222HnZmZkHxxzgLR94DnRBMl
b2UaH8Uvnhytp1HSLj5iebrGrs8lWj3rsJJX4MAH1x2DcoRFMr7077qVZ3U4YoppPEuYi2/V1Cmx
3Cb6arCez/Of0obmGd7gEL3Ga64cVhjrISRMw2QnJokSii/iddGTIfRPaS+KujHCWqmByHWXfRn/
pJTJH+f/c8LEsokVDQvgsZfScDpEJW/uPgxkPlh9Evqabj5D8zIbzzLUZCc67/t33iIUF9/4pQ2o
Ub7tSJqTsNKTC/z6rdeAGptF0js0nVvW2iQNjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4432)
`protect data_block
4JE9HKR1wipuC1UmH1Xeh+zOkwm0sVxuNfTQQWPAk/f/pFAA4Y5UnyoBcuWOjC+xU+ffM7/1rfvG
WzSxTbiA6nyYJA/5b1gsroTul8SGd5EYAUOFXY+8hHWUSRxip3yyKwspIodLbzX5ns2cnihy+H7v
N2hb0B/ujNOSUhpbO5bwghrO/BUvQ8dFgP9eqfGKmVvXvAr3nHwEH+tSA4mWNLaSZUGWEGzGwEFZ
nuD4dIKNm1FU34tNkga71Jqmk0tNDPlUb5Agtj2vnVGrxrg2YdbCqk/Tww2gIFHF5CYWMQkPXcFq
R+075U94sarVwQLrDkFNgUC/j3Zm3zApzhYca1xQsCcrTaUT68xcBkKduhvC32gfnwqZXzmddWB9
kAc9iTzZWxyXK2+ZdPtUoTOvOQzt+I0SYIYYpU6Gc6ajyfOUSvQv8150e2bY+B4z7t06KwZxrSBe
qQofEc8HTRW6J30tN/tJQMXaneHBEJP7JFlmBRmg/AGjBbMye/BVY/fcNnrldt13/+5mYzc/LVW3
JOUu2qbtdIXfOiE7+ZaNhrAq5qy9FpSBAMrV53GJMqakRgKHviuOJfBaaz2kRVH1CxdKin2RFqqi
RMGp6yVDghOkif7R4PrXaQb8SZOduPp6iG7u6kYtDICLrQSUVKjNCYrjM//zOdHQXAoTvTSEGrZ0
EmrnHTNMiIYjSnWy7cayxdVaHLuqKCvNu9ByPXchk7Rr6tiLlwdoGahuW04dfrB7objueTpXBJvM
82MwujdrwQdSpTz53sC+2ohdDwa1HicNhoZpvwsQVvmkwoYvqVXp5yx63KhmbpfwiYWayV9YMY7Y
jgJq0Z5pw7P+PvMsJB7sMeQ/tLWJttu+uCjsyh2Orv+icGqxwBeJH/C6wFV1KMqxNWRwY8oul0fb
dXPFOCEE1QMhdE/DaFUhy2ceI1t2EcMzIYLXrYr73foDTQFf4eAjlAKVgXJPHX5Q8c5+o8urAhLF
t6YzGPS2vDQw+/9V4Sfma61TKquWLrXGa0eUNeNsODVAj9F/GsCX68S7/i9xU2E/fLwIYKSQS9UJ
lxvkaPJqZ++MSj+fxFBF9BlLMG8RWLs0SD7GFWnr+M4kVodJkGGXYC4b+UR72awj356DcLLIYudn
Z5kZ9GG+Fj9sb4agctHLG2XHx9z+5g2x7uZfURsl3wwSqGFzMOt22Ny5R1L1pDqvussL2yEHMu/M
fH5sMGD+XDaMVnxqEEp2IukCn+FqdwiyeRPaQ72oAIN2/RM0BilKpaCb5rNHL+qBDwld8to30o5y
N+lM6Dtwkvyp9DD+08W4wLPrUxb02ejFvkgV6anCxsSlUVSPQHoyW0WHnqHsT00KKk3VENxo48NO
yAkjLr+LQ5IFFl6r3jT8i12cgUZ5j84F6WygkfT59sHPK5N+Gd1uBI7q/A/QlFyV0hslbVAdcA59
HicX/gHGqOdE/f1UdlIrMAvgg+a57ka0xwkyGJI3vqhHsKNTwUsEVf6vEKqN3/uoaVcgb00guHj8
cQlz0pdV0yTwQF0ZbE2uqd+j7poPkax5oP6pSHfMtV0TP6ltil9Y/qU5dudDfvfaNIpYEKni4e3W
i+WkfSpRxqq+aIQpHsQnSPVAQPKHXCaehdi4xd/EUwAFcB50rPqnnsKUhiEUR0j8iG/2Gaxt+hAa
7quJ3j0Z/PjIMKkiAqTu0S+q9FGUNhmMHfWngzMZm+Q+up5oO/ZRwEl+nXcJ7KOFeyKDSwmgsHqb
3Oat+WFQUHfGDr6qEQjNQRC3VtNuepwqYMpG0mUeBIWreSIBsJmtdv+F3nEqwhwV+OLR8r31HFyK
5KC+BUDMV8Aa05YXF3q7FENqhjEi9No+rl1U3CjkpclcLomZSJLsswTXqkldUbP/ATqmnEPJy3FG
UTR5e+sUPYBTJ2RrRKmF5Go8K6ijqpDjebc/Iysn8zWRkMfaHAS+XJ0WNCFsbFehghkPxLFMafxH
o4b2zZ/S8/LDqHggzi/EJQJJxhEdeCocHIaFgWAD47ZBjmE3hPGYT0dzbQVOaZocqS8mFU3G6dcN
ZjjtbsFezyqQALyECIQb4/t3fz1Z6Y7zFl+b/NUl1tzwUUNnFBNV/ypIlDN4EQNxDyS9uCGnUJ85
mNT+PoVQAIbfvTyIKNBfbg0f4xG1Jwz5SC3ZyOto+erhOSB/ez9J47EuvLiv7oPr3Q7PeYQAS0+3
LWgyiHS8eHSu+LTAK+jCrPPawW9sfToOpJDLrkiFi2r07BAB5VuE4SI2NHZwdyt3jy1zl/3ghrjZ
dS4qLfi4XAag32XNZ6qviSGEdedMnSRp9In/WrwlGNiz0kF2DrWIqARWaT15lRBG1/xTH3MjvTsg
JHf9NcymEMpwyturgafb+ZRRdBilNvwVgQBRvoM8eHZCqIS4WsGQ1B4yG79s7FpH+ciEqKUlrN08
9geSWY7M959Y/KQOuLVFoqTvd9Qtdq1nQpVquBVBk8+oS8TU4pOtSQXlkHGFqpRyJXP7OS+Gl6aM
K0a2c/ZLTUhVlivYI7wN9QDNokeLnNEgzhq4mMupaDi9dOPSfomTloB7JQVmz3r9S4ITfTDGj8tP
PNLmn4hLG7BglTkkHW7hmqk+oiujOTRd18SgnWIIuy320mQL6vjYkEcHmGKmF128Hc2CnkXrJ+3x
fmPsKgKrzCcvdjP/bZZFt7HusG9rT0jEi1T7iR2Vg+JQDXF5unV3lH1h7U8xbOJlZ/N/h+diYtBG
VxU6IGaBu1Rg10YDlDSYxf2x0Uqrp8MUQ0G3C5S1O//z0uuxOgp0XBv0S+hp/Jd2kbDGv341d5hL
Za9WebKeA+78/BwYBUoTLjZ+3b+gOwt/FcsY8sw0c856bv14uCQd3eK8IAsv35/v7qiLKwabhmkr
O0MSPJpbO0RBm4lhaEw5n/Kr7o/jXVt2/ZcPpYaIYvSVovwSSUdy7sie0kyjATwiLHIIORhMLEY5
R4vIdzz80bOU3iA3vcj0HlvfS+rk22W0wzsmDzhmKNhIpm6vNnI5lPkZ2Xt6KFHJDRb2wjR3ACA6
xSHIFzHFJASpRf9KP6eTkqwxiSBDO+f5XozGQ+BhtMxGXF25lZv6TQhUwSCXL55aZ+M65rmnDxKk
9hRy/3SJ57H73YnMMn0tfFEjhy1Bfp22B+XPWUZD5NNz80bIMGu11Hyz5/P88D86tGn5bv6Ah700
3AHuJ5KDoSYNSj5VZWbEk72mknS9Nd5OZWV5Cb2/mq1J0eIIZaPKm5c0ipAprWo6FaIWcYR9+rCj
KJDc2jlCTNSI4A9W1HfZxqxLheMow81M0R48oX7PwXLm2dL0rcwwKXbQu0PfiQDF8yyZIfVzkD0L
0CQ5YwOI6EUKJYiJ/jPoZ3WK55pBtV8GTeD9rkVX6F46JdFpeiQj4jJ7H20/jLndnKwGF3mLRX1E
JHPv0eme76N/9jtSrNa0psWHfpvzXzEZQfdGmUmsgHGI244uVwfAXY0MQXfi8JmY8hZpsmb2gt9z
+uFKlqpQd3Y4dDd5t/qA2+a8M3w0ihSVZqVbIkB54VEWJQIm4mcpwNZLts9BoSR5H+qKfclC0OB7
YeoVQ2QszVKvLXGRmFOXWndA2UlbfdrQd/QKjLIOKrKdDUSTvfGchkMKoWei2DDFznw6+j9tPksz
ecgM1mr685MOlih0yOWL7m5pGT/rxijNd8O0WVfbbVCI4oAYFhABtVs5J8pbWrRtPssGNssAF+hP
kMSJVAq7XKW1QxFDJgyxQh3hAOGM4P9zJ0eUG7+9McawVOuITntTVSVQ7oFVoF/pQSam4gTmPZ4G
nucTulQXWnKxSoswNm2Ijc9dsEXaJ85E4JVFKGVJV3dM7gIQztDsvoHYBHXmlR7mgxV2aofcASOg
HO8Jh41n4iWYfhmJir8jcXHg9KN8iX41w1g+XNx1ce4IaiADEarrp3+uuXtG7UT87FGb9dJqQAnS
b6RKA9u/31U6YDxFs67Y9ukKUVjKLKBeyT3SMDthNh3shWxJAUqn/p0G8RRVYxp8XixgsqWJF9pb
wy7dGtIpW9Xe9E7wJZH1+4lqLjUEscdTaMdvhSRmHTEV19a5QDpQBNz6iaCjqy+s0RVE5WIb/Jez
1Hx9u+wY6gny5qqXQRfgilmdTm+wDFCUCqDBFKTY0/Hvr1cmFvPqAJe0gEKdoEcy2ody6snoILFY
+mf/g4Eoem1mirhmmqK3Ftqj/M6hHSa31VI1M1K6eZjCbFr0aCLCiH553U5gK3NXKq3nutWXO174
U3twfMmlYqSyyI8AKXi1otdvM6rli3aM6ejFvNg6b4fCYwAfT1BJmdvWur1uWASM3r379t7T0UV3
lWuY+uBYeYdimLIcREa1JWvwnOUMUrblSwUZUvw4oKoiRV+tKp9wmVQnuBLhuARTlxtBJNEzgtzn
PP4PLta36itRvH/xlLVu+6eLlpIHuis9u7mppuy8otILXRP5DG7EGfxGzzrnhgYvtJ/0u6rldfYL
ODoP7dtBsKxRSONbheDmDhpwR/N1Q3GaeTSFSdP2OCwOhgrN4uVnYRPHpVqSRFOvGsC3e4q5A++5
iK47scXKJ86SaQb+s6nbgy92ZSRJ8xC5dGwYmZ615QyRbHF4xJeoH373r7WG6cEnYSgzVmBMivAq
5xsLYgUxMR8cxMjZX3ujjZlV7ZwZAVj58eEQGnXvrVTBCoQlpFZUlqQAlib3aeK74U5nsNtANT8V
AEyWMzC9PN8bnf7m3UNvkiAVbihmiaUGozkI8lXgxggUB2I8mdLzwhaJwpiCoqcIhSSiy+3bmjR+
4YaKUImveI25q/i7ipXCjek2ZfguibHhelr6C47So3Rc8nvIqtFwyAOW4z4BK/TFs/kTIi/NFJrh
3Fj5AMHM6efBP1dRcKjcJSbBLfw48PxlkMrHMMYnngQD/4NrKn/34HB/gqYEbufGluSt71K+n4DE
dTsaTlj4t7Ue3sfajiQCY44aTiXY4c/7Rux2DRwVcb2vdqMI9z1yGdrsIbWWH90mugx9250dORoD
8m6p0XG4KWkDtGdGnUuOQ1K2SJIQs+GxON9BzFOvDRJRC1Le6vrm/SH2S8r3vr17m7EM9Ud7vQWL
0aFyNBuKW27PVJKMNMon5YFTPu2TXG/95OMUXMtJGMFdwYhhTbStzKoqfQ7qTDBzYlBkomf7EB6U
1qVFXD4BQmVXj1+2/sJJZ6Qx6tNCuHfLvUJAqAbD04SNevZT9cLwXDPhZl6XvWWYiv15eXcm4nvh
+Zxk4GIvnT4CZKeF+mXYgeOjGjwoc2k/uRQhTzqj9U/agnsbBAokH/SGirfhJXt8qYiLKVGnVcRe
wSdlsvVjVs3PBuDu1stj53Tc31mOVNYoQaNUpMPgC7nDbp/OpmglMC1I55e/6Tllr6qaNcz9HaIb
y4eC5feiHWmrie512iucSCWHgsYHZiZyHzB3IwIM+F3/SSy9MB9X1yeyepYmLboCfnv0brimAaIX
AViclijlnzq/omRgyIPO25rzcTITiHkYAcn5RT6efIwN+e/CEfaDUZifjYTpt6iayIvTTRrtAZNG
Gk0B7KXepirmdp1NB4lhvthc+Mf7Gzo/KjIXtbbetvrp1jYn6qoPREdPJRnA9rrxogtYxG7jDMbq
NlkahNvKbs4lWNBTjXapSjOM0Vpz9u8Wkv1DPO+uVFuJN/OOqkR32ofXduUdZ2h+AiBCp77cHAnj
ikjLYp3havlS7Z46mlFCW3Lit+x7efpgYDOUGPfXb9lFVSR3RtP1IxoIeJiPk2G44co5mV61cKlI
UaedhEd1UipdKkmDy9u6wtv2cSeD7C2ZFuKD8J6CQzzFt4hAFkNFdi5L83fgbTHel7LyNS4c8ia5
k17IsT9DIzIE+NtJhlcoZfF7ZVVuIpJZn8VIl0m9xHxUxgoqQ8oTaTldLg==
`protect end_protected
