-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sQbcNjzS0yEATC+dc8Q4/zOejQgK0LAaoweeVQC/vIaYcWDzKUX8ZzVSB2tGCpfvpZrkphdiXJRy
JVpY706sUsvZ8UubK2eY4oNoY8UKkjM4yPn/cLhBGuccr6OR8eDgVtPKIVPd4/xm2ptPEfdE6bsf
wm418Oi1jRySRFqn+dB3qkCE+md5ty+LQxoZfHLeQ42lojuEBjDo5m0leVSwWmyg6LR+dyOBQTco
rVe4galyz/U/T6iY5C3J7h6SfCx5Ed3IldmmF4p0keDchS+i3repmQ/Ha/u+WA9K0z1AGW5VphVA
jbchDCWA9e2afbeIpS+NtcWgOt4EOOdoE8zGPw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25616)
`protect data_block
SzibNvPMa1ac9oEJjet2SJFBINWUzzljjn2JcYzgjfaQJ8AF811p/BrRSsttp5GDJGycVW7azyBf
N8IdROI3RyXxagWnfEHsUA7/zLdSF+wJsHX7iXZ4jq3sjxIIGAKEtXfepZ6rX5Dr1bXFhHMY6TqA
muQphkkrdrJBqC6ruxMktjG9wKvY8tjYDpdxJCqpaTnFEjgEsMuPa4gUiTiUPE0blCV0t0rXTMT7
nkHP7k8nOKzjxxJkFHdbadCPkh6K73msZ5V7jk4G4/L/CHWyl7SnfSjQgmdHIG7x8hUe1E0wQ0Vs
7K4Fi+twu7VlAZC8Nn4ed7eOCYP5zuMN24BM32+c0JPwJ3L5mNxegJTOL1twr699ba7Zsja0cat5
l7UA0EprYwRBgGSwisZPF27+64wqu8umAoTEXjK3DIXbzZTwTVevTxVdeeAmVSZ1v8PLBlKFFT3q
ID/MO/N0ndPzJggXGPEhdUtD9xdHFNhpEdFLRjixLR5o2mQxvYgeQLaWFSSrtuf4p43rILK1IBW1
gvqEfiGS/DJLSfGOq9IxkYne6nq5YX8HU/A2rU/XuxqBsNvNEled62JH8/XiPK+rrFgZnkA0fw0c
GkKyWbOMoki9I2KXMH/r33gDdFwdaovFE6fD7S6yfrKZ2vpzkgXJG6U7c/Dxaa3x0tTwJwzlRTds
KhC/E3xpe7A5LSOyPeKCAs6HKtZhEHthdpujQig71JSiQubEu3NKXxcLFxUzabqr10ZBmWfwaIy7
fgOn/tx0js3eh/9KNTqESUKN99nnMHioJLghNn98vmnJNJRRq7scs1xjekpd7zEnlDkhSNHFPn3M
278kGiRhW3xmnYeuMPtkyX6isy8z1P45rnnhNo27oBrVQUuQp+hpYFtl6DFIaXvOCLq7QCJl3+Qk
HbwePVYTvI1830rIHW6lgwqIVewMvGqukbF0wlFkt//zAYxRUeR45yYSdqOI7YW9ap4/DVxzJxhh
XKoUDRuPRRAViG8Lmjo9JttE1MnqZS/NfPaPMsg1wzWjq9p/A6jMJa37d5xcQ3X0szmTKrd8DZ77
8ZK/KE1zLuxtVhz41wZRVFRrOiv7bLCtJbRhTgNEHfpv3lCQeo+nI4ocmYDug6gm0bJCMBj+aMRK
s9IosT4O5AjoNCY/0kgBQDtm73bZKmPQQtWEo8QTRjRk84gQYlDg6lqZpokSz3pm8xEyDkiEMKKw
IWFTBPjsfSRwJgwWq7Idrf62Qp8Tbs9CcwQgaLUOI5trb0Hoqj1hbUezuIx6b0P9IoyXXg/uyIK8
QGrak8e9eXbmLWr/2ROlCk2OAaxuZoxgh/yQ8wSTqVVlBVSZuyfpVlxZGW0iZy7NUEBelyztQCRR
18TE6QybINL67nqd7VrhoLq8x05II9Qgyk2+dVw/DVdWYNzS6fpCSXE1Kc/ph/tWpi9n6CH0kg3u
zSdJQ8sdTEmBkhhDwCDXwndtVsVa2rk9R0zZX0g/tLojqnslFLqIURPw0L4Mz1iZ6Njb1bx/MBTG
eETIUzXmOFwIOYsPPGnz+Klqo+V8cyzUItjx2FeytFmqIsddkwqb+BplR3tbdxgT+WygtIwocC4b
lWzMinX/alE5bIj6jE7YIqjBBIatFIEVfYG/8+mwkbaUGnRQ2kOgjfJb81WPF2f1OiI6f+nldgu7
2fkOqLl20/el89AQL0afHGRT5RDZY7qt4yXvMU1Jzdn+0rCIrl4TLPz1dvksnUfQmYJ1I8fDruBe
Alqul8nkeFLm8KdysHtTvOU1IjRgiOe+ov82Bp3l7dySZqA53cQrTHkQXTZN4SbgtggZ/RlWIV/K
FtWJ+FX51TxgbFK38vwa4JORYiLQfHy35i8rqnDW1EfAIg4GD2veZy/HQgA81e0p+cCOXXQP8vXZ
YfMB69c2zZBlDxqzVeyFWdbW/8BezzYBlVoZTg+rNgAlXy3NppsWpL6VG88G0VYx+jxgj87lhuGL
fAGsowB6m0nD75NrZHFpFmQaXIm011Onl50+/Zk6B98lvmb1cYLYMmf9dkHaqjRjz5MT3PBKCtmy
eX+BM8BXX5muV24a4K+Duvux2FXLvf4ANqMfUKZZl45exrNsLShgxUAky5yE11/yQPHXSIiAPdGQ
kj3pjOdYzT+YDcvAN+GE/GTDsb/CiWAT2worsX6PriuJMXvw1RIbxVMJKg/o8/ljoU0VxTvy0ih1
NR9rrQEz6P1fhZdkTU00o31cwJrGqkTeENuagyhi9pWNQHZUjSt1vGgl8Jvh9MMSTjDtVHGN+e/k
WweJbG8o28Pyf8ecguNIBQYwNSbEgbOViIcWN1wJ/TZMG53QFL/83+XJcKibhw3opEFXOPM6JAPf
sCrTzs9YkmzU30lcHftSvmLzgj5Z4A2t9/B5+uDlcQs8+60TuE77OUMCReH5BLYRALiN0daHbym4
HOAdRX8MreXF1dwaVQRp5cKFTojcMk9a5es6eElByytpeO5cpK6xJLazqxg3wxMxahsgRCP6ZrQo
1aRbU546da79YQUaavMOmIqxA5bpixLVbl54LCFeYrniCuD+yb0XsTLqQG5oguUUWuW7DDXlrKQ1
onGHEqAADNNs3iVj6rzwLRQtusEwzEx6Pb/wSdWdIFI2XW67n7QRri0rs4Z55eKqTOUERU9x0zkX
g2XnDYH6wKNtrVElWmKC5hQVwoJcIMVQsm2JCwwU14xNnK8LXQMSg8DaKzOyDCHxXBCDLGLy0sQ8
DTaXR+iCucibP221x9s0MXjXdJDZxfVXipf/Vwndz8odQ3wFl6Ob4QSaxn6CzcwuU/VdJSrsEakP
U6QUfC741XFzP3DceiVim1O2S7u2XMnlcJON/dC1CyQjL7h5FoMZlxVj83OH9+1cpjZXO4Pz7pe1
C9unLrFRYXhVSkSX87dF8kj2Z9Lk59dvpS13Z3sLVlLAo+/Z5zQd8TmJlOQoPV2OX2/JEUgyhOYD
BUczgSDCfg3Oq9JW0Ee7mJZ1MfiRlBlzGp8oAmFKdMg6PEl6qc2mM/lcV7Mb6B3bUdchquWgfIum
jvmVy41HeO7oak5hEtrXIKN3WOu2EBVl3QqvCnPIZj4jyMiTxhcUY/pokI3G5JUDqtPMNqAA6E7r
fIgdaZSiesawHKGaLwDuklr7y9eItBFiTWttdQ5LrilThWP9r+RAUGGO3zMnlk1E+2ZR2e/Sdh75
gRQgSGI14847XmgG5vqaphdRpa1sFQ8UO1g+TtpgnHp6YqOOlr5xZO4H7+P0hmvpVI2kblrA54RB
zLDIkpJpZHgeNK1L4XQIQXnLlxxpJgiunaC6nTsZ0lq4mjKPEw/Zb/XOfrgRn2ayshA0ogu+sOtI
HtFQzYNheh8OFC+MvmP/Ju/2zD0hBhS1f/VsgmVddnZ1EmFHrIeba2jHRujI30vtjN0yRx7R2M4c
6pEjTKT2yIr2g64J8xvHC5czgy6IyqLK+5h4NReOyXhEqXiy7ZkVtIYJOQjJdwdqAWvBUyGXqMr+
5q2JNb/EbIooaWxFmYb1TXRQGATtvahQ0fIJospXyeIDpxpNlPnYhoJbdTYo097sYgzTD49r4EYw
3Z+NEw5Psd5d1fQDK0HjIzKGNngsfjQV2ReVgUOGecGJbPBtsBH4PvT7QXhDXzuMLphjYq4e+zP6
emSG0GsOrZEM7N8UiLPQOR4QKv7lQjHF7w+MJLb7VlR+wVfCsoeajBxvGN7LkYvQnrHi0ivRhpOA
OHZoUkLkjtVZT2PCct8uPscjZexOclQtxFwcPRT2DQlfdLqqt+ET18+V9UEGGCVlQiw+LN6B2ivk
KuWStRvZHFLON/y/A18IodGxUSBzpdmTZUn1IP3FuUAIN2NFuF+LoUeyTLeglTc6nX0a+WZbRXte
I+vZ8XHvdy0IetOTT6n5tZkl59uGt40Sgo1FaQwbtPzj7HOmj2VXHkFEBH17MpLcXfWW9YHCtxUJ
rjSY3EQxcf0cfRqM9WXHB5su/+uU5AA6+Hgi3hd3/ycSKLkxFVxpjB9165boReFHsYyiXFLTafYL
TQS3eEX3DaQpQRD/9kciL0Yi52YtdiMjjxfeRQZYoLg6QZfHyFeE4+GfZ9jfCa21L9h7vNQsE00l
N+8Hk2nVCyueVJ5/04r/FBY1SGOKD3bhe1HL4QIEFM+E7tBLsgSBZn7fMSpyvVj40murExQLlV3o
D/kkhSTVM0TMjczt0iiq/OcUthqoM6mYXimtG3OwJFtc3kJ840Vqlf6SqpTUdQmGjpbAibngAVUf
HyOSNxB6RC0Bf4o8HpJt+OCU4ycxZsgfAG1/KrKG1dcqEe9zm3wmccBz+O1TDw6OblXN0CjmjUym
QiGp+msBlDIQ/LxOgdxnTUWT9RwT4DbuSvlba1cj+OfkGiLGXr1dkbt5LbfaSSoly81Xw61PDDoM
wnizYMbuO0rUlteBLyEyWWMEJGSiU0eOEpVJrskbNiYbDzIY2srprJQhEZ03LjmMFdDYASQfsvpm
XS1ssJPBJehx8KtWQtIloubIL38IAbYB8+VK9LUrw8Ocz5jakJkSNWBuOCO0wm5lrB2FsyUGZuDQ
qVeq6uw1BhEH8N8xG7uTiQ2EGXu+8USKB6W0U5j9pGc8V+oBtg4mlBxUH90vBSo62EGChwtsHUr4
lPZPBB6sfBJgvpg7EU4am5LSJCL40VvSf/AvKmaM9LbsEr+PtL8CLVdagwo6GikzN5bBwUjoT7Su
U09BWFYlO1AmHboPTXtHfFPBJAGAv1aaiiEqH7CMpvP7G9J5pFE3S8rMVdQeIUEWk0xtat4X3FPC
m5GtpDqbn31TfZT1OjdFoU+boSJZSCFgvxkJJHvKcLVjt2uNu6wVJlhuF/qe3k/y0+O/cXriz4LJ
Unbw6P1W/mfvLlCgY6pNY54h9MrIFGLCA0cajZpQFlKvp40AFOFy17IvwGiDg6AbYYGscyprLM+1
8eefn4jdAaIuAb7aDKLEfkFyDVaFGQvtB/FJSPBmYfc8d4bFcKfdA2dGVIM6wSVnkJyDjQKv4dFP
FsoCnKfG42DmvC9z5PgaHX9ncXrFg58+MRWkjs6C5lHH2TtYFISHTuso0x475To/BJ4f/K5w5IGX
zkg2wJDztdbKcxCXkFG+qssiH3DRF2KjqVct+k3PR78J/4zSy/HEJQmbR7sSlZm6BA8ZsU7RPtS/
xL0w3dQWdvsW2u7QyKx+vWPHqlVAjBP9LwYtuvRYge8f+6Djbds+c+cjrViFwaHcqJ457wqQT5Y2
TvdfzPnaVsdUZOv1detE/9E/mRjg++jPUVsyEYuD3m/SuqNkSWcQ46vhcTCiqnpxOHT+xDWGqLQV
B8By8bh4YvsDmUMUpjrBa80U3TV6hmm12iXn451ZnR7RzYlcqc0BX7ngVVVklNymFPC6QQyHuM7i
LRpuK5Dhax/JwhU7b2boEJvI2LQc4PQns5UGJMwvcXQJYzgQzMiWDfSSmSeOBMM4iodIAs0+CxnC
ySlNN0VTdVuicFsrLnvklLZfxhdbJC1vnvpRvwxCOMjAjBWpnF3CUeKytyLlVNI0Lm5WIAkL0QfE
wOpniSqIRa0ujTa8dCoLJTsm+tgrCNOQ/bQRvSHIYfxWh2BVyBLxq8qFXtFWxHT5YXlqc3dTH7LN
gBXu3V2o5NQPdVbCEE3gAD9tGyifLiN6uDciOPKtJARE7826+eE9DDooyIUE4HLaepWRS73sUMr7
Hk3JvGGJ2ssAhelr+Gso0kFAgkNR2+34zFbvFcVhcuaodBzgIVplveTHeIDczakAC46PqrEBtJSj
YGALz3r8gDz3Kn4izu4MUmvy4KpZQ+67zei5cYsAYi9X3yMFeaOacI4/MHJ6iFjYUV22bvckZXZj
Oz4TpfnWP47J4WOvDMW7ZhFVuI9YW16+DtC/hRqaUHaU8oEP57fEl3U1fEBPjmGGCjaJU3XE/wkI
cOq2W2agbsY2nNGTADV+NdtBseitXK1uXPiQMGunEGO4Iu66d/hnvq3a9BJwZNAU9TVFBzg97QaL
WXz6R5RUViK8paxaqN66W+9y3K7cIH0BmllKjmAcUXMHfzv8tP6SdNUQJlVx4HfMyIRKXW78/Zca
OaVelcHt2zcQJ4tw0DnhaCnPT8rELWDZDiBlCwx7gEQzNp66WDrVDK5Zv8IHy7AoFJr1zclwYx90
/uahwaWc2R68L6k4kv+Cop2HlO/2Kj9h7iGJbh7KyZp2IaTHvGzGU5FIxkQ+ekYVXXQOgkFYviYa
wMC88it4t24ShRWWNJMyUNI6AwRpxZR6kEhRjW//L5+NrG4ZVuMBKKeNPYpZZXTvVNq4bSNTzJl0
E5+GjxMnU3qwa2LNqTyF9BfDudl7TExCW1vJgLZq5GQnJ+ZnYmsSaD0LMdmPJIGGmh5rLjkpWaXN
HpjJunTINPmg+AuR2ZiA41GHSsU7raFaz34CpuiPypfYSZOiIUgnMTgojTdfQoi+mhiGt6okvL6r
VdD0tahvLfuldYR1bywW+Ivbk5sFTSVbPX5pojoD5Ua3l1bR9NLb6j1Dhq2okufNeWgmWt74HY/t
Je0NGK0Smi4LcvTxU8bqb8+JWuZoyO2E9W4+oubS8WvCLZjNaSUH3Z2AwPO+TogbFMFLckDhQ4lO
AafXSlQZU65sCJxLv4Ybtak1ZKk9B/RSD8hVVj8oBOr7KEVvhdoIJla1v7NuYzwtOQBGppbwimAh
1nJLsDn1ma+p9q8sdNfGTxfuOKFUdP1B9ftC+DLZQIlid9sfApQRaLhDBhNqg0He5vcldsu/qD9M
wY1qh5EdJwiJEvXNDqfhAaHWXrp7Cc4IBEvZSExnk7KoVPkqJoZMi3dmP4VhPCAIC7o4yivo949V
xGROkZI6PUNQKCN4C1M7KM7oAfwzSYZ7/RJwgtvwfa6zuqWc6hw94fOBPZd/7d+8KuQH73bfrgQa
Yyv286dKbEgS19nQ8Ct3OJvc5fIwzlQnUD+mXjZ1muiHrYOhettHJaqJqtUkRpfT+/l0g7Js2lnc
Z54z291yQ0lql9o2or03u7aFnT9/ncziyXi9aCY6QQsa9MhWnlip2iTyhlOhZ1nIThzGqj3nq8Gr
mSOWA0VFoJMQEdsdmiIuYtfQwRsiKaVxN3cO/tnmvwzYQ6S87Fw7MU1NomcGzSJbImlhqv1gOmsU
M/dnGArrLBCHaZz7MD5up+w/Qqaq0ASLgCop5JSTKfeOxM2dSByKQBKyNiNRfmcOS9Hygr3mwLst
7lg6BfYoaL6Fwk/vgI4utUcgsq8DmkHJVzoMwFA8M0eCtC0OgtJK92QlmdaHGxuXR3b5v5KQWVlR
QGTmRBBB1UUlQs3Z2plWpcP2ePdAyXa7V9xftF9xvlv8N5nnHDvXjuctWBI/Q0yS/x2FTcC75lo8
2TIoE/n0JsKlUTgJ5mFXcOoBpUymHQhai30Q+zP8OpAcjI9CjjTs0ql/zyZdXwjxETD7B+aXA6KH
wJUpmAopfQfizhfCevdgdMF6XAQdHrWiEeWtozwfZ6WigwtxNyKh/YsY8cOdXNjPvO/Zs+hAsqaE
iAagWc9j9jY+ktPKsvoGReHB5w1C3/Ca0YBzLTWAeFlOEe6AYnj3NkOIkztYUNgK25o3WJR0XKne
SH7wkRana5cYosU3WjuU+oOsfAfbAAl3Dwq5eL8sIcikl3kt0prnREXFI6VedKNpLNiMS/uSDdCA
xQjDkjR8S8T83uIyJjXwO4yzWZUjBAnP8XGkGs6xpDUoT4tacwbMZMP4pIE23TtK/uBfqDhdzvqo
zbpl95NJBMr1QFuGdghO8rg9Hn//MkJiPUE9EMhWK408Z18Lz48UK+9aTJLyoiWAty90ftXT230m
v2wHpNRjzRXg2TsAc/Wxx5QvqPyHwIu5RVPIALzjRNttiou/DnYsCZ0qusS/c98hVQYFM6qNxf0E
XEGePmokMis9EdYybiBLjRmKVLF9A79/sf3NchQKi6PrDkjDxpu2pq0nBn7GF7BslkDy4TKhoXqj
x4cSEcxycMfDMKEOirmiYzMeSIzAdWPwpY4XIBS+zAddw8XSyF1YTk3Dm8ZMJG3Y7TvttgRYhOiD
HFaAdhiu1USfZtPS7ebO8wdPj0pcK+GQP0QPB86IGntRqXFp4srRWuBma0ZCdAZXmbtc98qyohSf
oNJjwcBS32ucwlokebW059VQfwR5XNA46ke8TuJlX5blx0+Huw2szTkqy0qv5W7MKOvPHfSClF8q
0+CIi/rKBFmRTy0fo1y7UqfT64JKvkUlwGkxuUHhu3IuaXadaFOhhCwfVTWuV0rLHTxJ39mZqL0F
kIH3BxTISypJ8mjTnRe+zjNUVpkRwbZ8aDAlOlXF5S8mI5LpBF4HqoEnTbic5VbHX3qM3rC5lZ/5
xDvI6D9TO0ppGuFcCdzT+tnTb39Nb/Cgax/bwFxcHKcJbnkHKs7x6551XMAreTM9B8aYYUGe/RKh
qsCK4OqGGnUti+hqjlLxr6sOcOnYIdUa8q1tBGmEP/AJ+buUsR2eanmXTr9GfM7zV+BgmLHGGbhT
wZUuVvPXEFqUOZrRoSnYxTAAdEaVbtW8Busxf33Jwi4t9CgTVckM85teP3PnKTZcJmsCq6BMrCgS
WDL8k19LHHajMvabE4dMeYWhZIl5UJc9g4nY8m51tIQOj/uyBIWNPEpVVDYm/N1/O4Gc8qyNjdAo
+HsWl92HW9geDDelSlUr1kV9tI/ffHIvGF0pVJ22b0WGJ2IntFLUtLxXv/Z7SdhYuU+gTZEoqMDy
HstLOu+aPZPZoUCuqkYlSYgg9DLjBUWK2vbLER1cxzEczizM39F1XK8Fu26ZEiHp7YUCYbzty+V2
GUgqKfJEO78rhtgaZR2ekxz4xX6X78APb+MDwVXeSgMIyMUYiBXXIQnotXMMf1/ZRemhuYGRVVkJ
I7JzKhMkxlbZFMh7/dP2oG+OyK4kbdLr7iV8cFY+YKOFrFFoDuO3P9H1BTIfswWhGXCmHoy1R4Hc
5eH6v3f/9URfAnilCEIOzeLs+dxnxGAmhhzFg7W5hcsDUzY/BSBoY5G7s3Fv/PJ5Ynv2rsayeC7T
YSApAR18D/IVPS0IoPvHNDRpU4EmGC4ny4JrsNSCV9B23bfe3+8qHiiBhEbWSt3TH/dvJfswotEh
pEHySYIRHfPCOlX9gdmfKCyTvq5nnFitwYdr5K8brhlTOnGmVzYpSsiltBItMKFKs6V4iF4ntJwQ
IKb1B/72U6LpuBH5HRxdskj+BDpAo37+xs66JC6wxDnnuMW9RH9Nz4D/ZLgIwJG+/AKcADGXJjjM
xSmGhPg/JX6fAzhGasvPms7vFivnpOR8txF0NOMZ7aI61l5VtDrwq0cmD6Fteyni7mdslIhcWxgd
Nmy+Wbp2OpKUe7o6wEaQJbOmo++i1mWhdAnIm8pYGpFgkQY2EbO01+KyH0pvvMBlPOqPCWKIlJJw
LEuTcRS0XCYVMfc3MBuuarPhT81b/rSOKW25pdj9FJr+d9XuSZKIgtDE717hPlLN0zzEvJO0UOZE
K0TT94bSuCR9Ak6IsfbnTmDFzKEUtMYi5BCa+qWGPefA8idI47Kx0IvK0Yt4qrKpkrle/1h8ZhdV
JVoezJkx7Y8hNsOOx0BukVg1o+TL+OEBQhw7XBNB2fVtyxlTVd6KEEeimQPhMdUilt9/T9gcMGFl
zT3rx5iPC+PhAcoBcc1w9kyEvSZ8R+A4/iJEpbtJAwBFXWuhm9URDhm+muqqoI7XuIefhK9+Cjye
K9PCLn4BzG2lUXZvXEu8RZIkTxVwZlnnLyJ6ZvBuWU9BT4QCQRaJ8iD6SWng1BiqgPJAY9HyB8ha
59GeWL1taWoHoBb3luUugBJknZelq0VgVn+7RMUEtZ6vmRI4ORp28jayrIe7j98S9m7GdoPp0I/R
wROb4haEqWBxXH9YlTXHi5evBz8CIs0rbG62t3g/lkCDiJpHXJH9e/rB7PkWgAiOXlsUjoNJlcHt
UWp0syCvQDUSka8rkjLl9U+jbzahmPRGzE3gsBq/nnzqM+/I741sjGXTPor0c2j5CFC2absRN/K8
Xqh6qAU+1cmUL74Q+dNaQvN301ZCp8LR1GvKEKo9zQQGahkRBG0f7eXcYVrzxDXhlmbsGmalMe0t
oq/zj2ZWjZ2t2fIDubokAyLJQGvXSf31HypRBHGTaPyyKDABcfPXRpdQu0k7r/9KuS9rj+23HCEd
ZGoRoh8QbLKiN8H9bHe/J1LdXTM0OJW9jqQg+QZKDLLKJXwema+hTd1QXeKfoVG6lleOhmpFKYi8
x6KUpCh/wSwJkbKHHHiKLaHfWgaxBWPzY3PuCDD90bY9tCCw0uNUDoHDOEgROyOHUd5eMMLFtDCN
GPcK78J2lLtCCv5VANi/NqgzPNO0YuFF8Sstb3AwD2CWC9Q0G7NnRu/d4l1wPL162T8ku1HusO/M
vBN7AE+sORUQPsGDFo0tv5NI65Xsbfc9V/UvW2F5DVjnc35TAtQ2n7szmiQS///BAJGA6wd1BHNt
TAHXvj/6j76zYWU+zn61MwfSsq4DVSlHTtBObYdvA6wGKyEjOT+rGaq1S9YcxbZ4jFJ5bF4Br6Su
8x4CYf4ibJZdGtfllA60eGlkf6uWsojMHJ6mD3+nXXnKZhTfpNMBpMAuRbiljva+48GeaycKZdpt
m45OtsbXzxVJTq8tqfOMrN+LRWCUWw2xYmNbjYhuOfPz6Vwr2LugttDA/Fj+YHU+4J4hTHoYCy5E
s98Q+SzwLAR5PmvX7+ev1AjD0mPJx7FqD6j3VZbLUJQBifu6+KfmKDBXff3Q12wVjIysDshCZjI6
B5cYLb9kjpjO9Apeyb5u3BDGHXwGNhSgJ32I79m8UR34QzqR4zwq5/O2eIKxDLlwwc6/cP/W89oo
8vFVeN4OyiHRUCAljpa4suF14AQXXM5HYL4RbduEVjpxbVSkvBictlLBxjuSvJzZPmw+NzUHH5Jj
8e98iiVIisD/tvAZqtBldVLHTXR+6CFYTpJ+UAAwLogelUd5dtnsMaDc72tBZD0a0VHE7UQ3jEhO
pay/WOx+JUIKQwW7slnvI8DKTJXod3P5HObyQoA3dTyYGCzpvr1okiWoRqVUeRVRmlgh5EkbqhFt
b9aHQnW0w0HqAD6Ueht8s/OpoMnwtjFhZevxnppkHrut12XAlIYSK6qaqBKn8DU1JIwmCZxq0gEY
UAFU0qVKSStwsU6AO2TOVzljuUjXu6dkuUZ1bMuFl8kBqWmxUPEoL0M5AWRNVoKG39dfydb9D2Oq
8105C2a/Y7Ibvwxab+2rz4IfQbRYLgXOew4PSDzBytv/Coa4du2FRFBxor4/Kux5fnTh34/lbW+p
QyxU7p4JfJtFbqczs4kwTDcmGAry1eLkdSyBcFOGTwx0fEy+rTteJ6rUcBNutUotquOyVhO20Es4
uHKV+ZkRqFW2iUltfZtLj3zjiDD7GW2jX4fVvsDf36++ckb4nxbvlRivdAqxR5LQbieF95mrTv5N
hjJhqizetE0mUGRFjJ1vCcdBb+fid7f8TkM345NoLZddRkIefz+HCQm9rvhrtQqWDVQX3YLroGWE
lTJF5aY2NzuVf3vs5LZLE1JMq2BTT4vPe9jT5M5O4NgG/Ymlz/KAkD5cVm8OEhvLvIaOODCkLwpq
m3Inv8Wcky2eEHKengLtXnmo0nA4zXWh5F8qlJrwLyoeDYG/AYajf2q5HHt3q3IXZ/UX8oxjgUEs
tBlOMznZg4CA8aUcPE262eOp0VL6K8T3peSvcaBD1HNND2T6eaGm5+6UsrA6NTQ6WXjHDWfu4kw+
Cl7KFYzRYzPhQl4pODL7ahqexpJyHweH9ve35ArPNmCG30hT7ZT9K4HJjktwC12pAxWeY+EOy7JE
fRjSoLajl0fYJg8JWBWcCIizLytx0DM11I7rejsKg40Yurto9cu7QYSXZVOVFv3gaaF1ot/pKV4+
Q5vhsDiHoXtpxl2HrYvq5x5olFqly6X+aiQwSHwtQ+0Lp89KW0J3QnLgkIZkfgu/HyKc/W51SATv
Bjb1baNrYp5kCz+1+RMosv3Xyv6dmtq4lwCVzzcK2RevEqpTwGhSk2w/KeFwiwi+Kb7qqVvu30N9
vRzZfR3G50POcphU0LaqXotnfCH1WBOCWW6uyPXderyWvAynyzvCp/ZTGthrAkC6enWwI62O5Loe
/W6mDuoNAw6RojuwLCqXbdNerda+tlTNw7UlLazO6PyaLBCaw3A0xmQh63n0Vjdbx6LCLE416HSC
YH8MhvBXMDDgXlhtG/G/4wZAWxLJG+M3uZtqDQVa6lLy03b2Cev9SHUaux5k9+IMnhm0meuIiPW9
wD/aBo7kq68h7b4Ym99u2z6T2WFX8bndwwbPKjmIpOm0l/GS6efOZxfs8gwGTe5fJlUf8lD7nVRa
gMRY7bHQvIrwU3Z2TD7piOptUrNBeeg/0DwfAO38SsyH2R6LAyTx0hcxwO682gTyH7Dy2w7nYZ8U
yfSGrdAAn5PWrWEKkD4d3HmM37qZwbkBcQ7oS8NseQUc2NIxovubhxqgdKEWWtQ5wBxvKb6FTOSC
n7GVhiuVBfhKs6QWKkuHEbfjxh3Mpt+CDTX7DAIi3EZdlFnNFPLzC2NN+hUuVoVQK2kO/KZ55PvW
L/uEMAd/tmKenOzQwILpnv9tL4p+uqSbwnXBrtOAhZUplxA/cE1KbCYBo86ooSpoQCgWfOXIGfLx
AJdEpwciAqfiA7y/L/wub99Gkkt4/woZ8Jzk+v28A6tmSj/9zqXKhOTY4Dog5UDh86IymCz4rUrz
WT+U0qq6RpHPv0MGrLzTwL+tLyMX8rkFx1OIasNgHh7lAL0WOgtLcJwyMLYJ+KZBvp/DLnSRPtTa
uckm4kZO2kK9rVnE6yV2lOo8GIElG8S2qQwSgUYvroOq1NY9pMmxQPG5SHH4ZGrQ82ma7woAN+Rs
5iRj70M9Y+rGUavuomt0KDHBZWC/49EWoLWbxQYFWEhyp+9wEjyIj4BaPQ1yhdLCFQz4UQtxAR2z
EKzbmyBW/50uC2TopthvbBV5Mfjw8G4fmzsMCuitpSibGr2M4mQLiMW5G/KM5bW+dPaY7vyPRkk6
iJBTCENTx1oo9tMVCoOmsR2kmT6N0BAEeFabMkkO1Tv6jKMNQ9Y4YhEayShBshrvpuziQ7XL/rrv
IlOJw+WRGGi3YIGLmadJBNPERQi0Zq0DC0gqXqCFkU7cUjgUtjwuBY0PgOvwd0nDkENTA1bMbYGV
3jzkgWJGveHowfNi33d/K4mPie4eKeZomH24X7Y3QwpAHaxXPXIfBzVwYotQdniTF2mT/pcX6cMQ
0EjxRayo0PkpcxhequM0aygKtzQPa/1DI7gYQT5m8UzKBqKtthDvOLnpryKMKpzMimFTp5wrACQ7
SKvBvz5BdogmHMYMpHdWktHI0ulawXvJLXQbVNCLfIOUsj6shlmRF0GcfBCd2NUl5W4X41WOmB8i
HQiYJYPwHzNaNpyJdV8hQGqCKGl4ncjWRGIcWAoq9zmkeQWNORUigZBuGgW1EsVNYHQdLLHUApRO
/vnfdPiMaDn3oAudEEHx8Vs9XaoKP3RrtUW6JF07gD6DTEpTUJqUFPWhXfRLO6rrF3WLKLAeYOBU
umWANgWcda/HirgSMTfjxGOhgxhlbqfG3ZgEh4EcAjIS0R63qheIF/8wJflRU7T4oThNY9JqY91u
vLR0ftDVxmQ4I4k3yOZDKMfzMA9hiFcStgVM+fCLgwmcIXqmLDU0ZAglntoAfaPFmM/q1uGXmb1v
67TQlZPcXNBsr/K/V7U/gZmAZ73yB6ISXJw9tu1ghEBxkq+DH+sr0QLD3oDVh4f/QvlALx9TI3x7
9JPhhdL7cC+XHPwHOc+5AP5xe773Od2r9F5WK5+CtELlvAkZddKiaNWizTWff+R1G6s4KDYREBgW
dd3xRYzGqyw383VWlituoeIYK1ICOaVENuV+K+XItab02AKxbUPilqFQ6XXxw4jEjSlV+22z+72C
kJdPwcBg6kBFitAVOWb1M1FIGxkG2CoLaamLt2EkPxdheeDQM61tGCwUngHuW8cXnFpZf1/dTfKb
xTqNhjNl1BAnIxL2RYQvi0NfbCsW4n6QR2voOpXopJ7hQBkJbrtwzpdCRLEVk0+czRUzwZmw2Y9k
h9M8PLHR8lBBrFBNJejMBzxI4zd4C8VDXVbXcwpzd29gsThhySI7+ZCmqCROA4Fo6Vts2rk/VHhz
s43EvXKdtdSfmJ0RlktQ+m8PX751z/arG/xU0mXwV6vXCY8VPPKsjKtDzA3EAiBc3xezHPqF5izm
OCJ5qVIVV2F3iJzI82QHECBJsQXHO4aOjN9hApcXHYUhDLCQkr7z0BxB0IcMeqeuHUQ5erLc8BM9
FpOCYnvIdwuxTSDNSHpI20BOD/ToyV6P+zTRaqHa3l/Rb6cdCh93T6mbbDrbBTD0SDUUbbcB3UR5
UIRd5XXYcWJcOadG7HnPrezikdkSVMsGBRujGIH7H3rgpwge1fCPBP/NYgyk5VAcLY7zW/01v8Wj
Po/9mKQ8nXvj+S6R1BZjbjIafxASdWz1FNWJm7fhKOcIKEBrrnapQDc7tbwPAl6BpBsNf0RugS58
1UIgZzykn7guHby2CjMk0F+UQHPyVJzcg5p9M+yTCLLC1RdApWKu8GhndSNB9kkTGA8tCO9BGcLN
bAKq6WAV8tD4wgfN/OmfYg1JjX3ALGR5+oYXHtF+FezIkgEwjkzhzKB3k80gFruSWIxjhJXRWij3
JC9N8g+HB6EGOAltEdVu44nMBs14ASKKaKQB6wO3id3++xlrpxA8Jwoh8sVdG7A9D43XzMdGrBgX
3/fA3Zg+1WbqXy+7ERI9Z7gf3d8i1In8gopEDC70xRJJzVm+cNxaw4aEKCF0RHwSJ5x16I9yXF2q
GAbt3XOB/AMoo8pEV6LpPNwrt5K98CHC5Oj+8Kip0utaltJ545S7G1WzN5d8r7VJtchRHGtRWjG/
7r3C8Pf46hkM960EIFTxH+ZLhSHqlCCcIGw4RVlx23LicV4PYkH2VD8QezyHWHDWl9PB5HZ2mI2h
FQcv8MJvZJ8qDgkAotQw3aEWd62tUevJKz4/dC7oUFrSaqDqjnGuzrGht0kIFWsEylY0LONypGdj
qAOoBL/gmvjSg/sjhgudguqLx/xv1s58wWSLdyyzjUunSc0Fb81ybLMX2zStpUKKocwA+lxpbhon
VIKeQN8e6vwSxLR0FZ0YBano13tAGoHzGiT4Ww26vZclGtIo6THhneO4rxiW9fPw85ifUOFmkEzk
3fji2wuECwfevz2O106oWEgCQegVsvVxHw01Mg6j5gmxpj9R8uh55EUMEfLMHHNzu5S4sPCU6Tnb
WO7dy4GVc1RCP9sBKEvJbYslobJ3fTFqgLyXmhqu+qYEIJQEpuoYSBOPaF3rn2Y7mQUtPcTxqwI4
eLWe0PAeTkiXtEPE0gKK4Jd/n84Aq6EQWUyePPUDtsFi5i2JedN0sIkDsuJs8ohZmqAQZQJ0z+uQ
zZRjxoZMSOItreLCJBQ/s07ktSakXsTcieik+JUVytsdlKYJ9Sbfj/e7NV45+ZtBgqSfJMLUtKPr
85FOPQSX5gTQE8V3u6xcgRtbEkeJX8nzQingSRt4eEoL4GdSFPnfbA1dkkkpQrHFcCXHq6Cp2xEP
SWrimkduldo8VjpkKJ9JmP5lHTQ4tEZDtN82JyNL3+TZVYDmjTsadQRVlAhPEd8PJ+87BlY5+Vcf
Z68yywFfunZSTfYtTm6YZz4qAy4H8M6CrePb5gsgvWI7Ojs75F508wovmHE6CFoQrTVX8uGTAW3t
cL09xnc9Z3ZaaegK6uucedRHXLUUOF02KxGyywooiF5q5ETIJT+JcrOnfxYfMWcWA0spGqs22qMf
QZu1/oX9hhOflHtJQO20LED+iUOM8UOKoCz2OHx2nw0a8Glz2X4vCJ/SAHPY2UH3LsPvojD0Dhf5
/NN4nST8bivRQXOwKMqMHwEQA7AQy2qmRjrO/ZalgX7Qg32XdOVCVmwkIAplTHFEg3K05S+18c0U
0f3HkNDt2BIQZxN8PRtYksrDSP+abxxT5pPKE88wSdwh1ucVlYNvqne+I0iVdFwrrWX9cYeQ3n32
mriTtMPCG/mOtg6Rt69U+yZ415gYb2/vugKw6VW3p9S345JuOJLx0Dhf+8+uVOCLnJQV7Qylb49c
1cBfsZCOIMWIQSRUKU/3CRm8EKjoLRH6CiYewZb60QGFUCB2laJy7+DuyJX1KueIQuaWkMLfb3Bh
SCWGMDetxfYcuFfD2c/3Zfq+LiQ2Zw4QtV8fMUpj26QKiQz3xGvomJqF90/7WxW9xxtyHCjggqEc
ofwHvwjskncTUOb7OJvdBrrQcdzKF0/oqtAUSZGsTHGLapfpdrgbe5ZymouXsZcu65G1EgSqhx87
s+33nEQufZ1qgriKiSfjmiOqWsDZ61uB2tGT0bToOkAK8WkAH1exKrqasatX5BiWZjakc2MakASz
D2q1r9xMzCtqP4u9F786fYMPp2nA0xgzbhh+qNROf46I/C7UYwU/u+L/FRP/pw+Y81a1IEbE5UpS
IadKXKGJ3pwUVWhEslkLUKwB8oGw/K7a8BvBf7Upsn1CL9SEQl8mcqQKAM1AYllpDekScwDsYQRx
lVWcKjdhQ9x2kqDg4fhkfc51u0/Fws1qxPOPSLVAOcuBldBGZJIRKB+iQ9/ah+qpf+V1kHGy4QSE
bMENwPHhIQSZ7r339jgCZBoF/ITvYHvDwLs3ddtM62TRcp8kcgfDZJoQiD2IfjYiZr0WsmXiO4X+
XFaInXL3fqnX9/CtYh8wsiN+5cq4jfj6/bq1/2s/0iMPUNaljSaRmguGUHwYlxqJYEwJXA7LY0bJ
SGGG7EG+pntLDeuQC03W10ziJqsTlLUu1/A5iBAh7td98/2geARv4CHV4jxIs4gsafDlk6AH69TR
R9p4AEFMC7/NYvMAiM03S1/NNRTVF4xOf9H7fJdmchQD9M61UgjCoZbG1sio816dYLiF1nE+YAxN
ezqG2niFo6ZMobiD1k/znfLynoMzNt9qtmPGaVlv8zycEy5xn7iV6CKRkB9P2xA5gn9fPU6m0Wz7
sSKSDRAXeYhicreuxfs8KpD+y7H6C95QmFD/8hpKcr9bQFxqzjYqXb1Jn/I4vq4YCP3xlmIh3sWe
IncyhIwITsfjAk1Co/m+Zq576vt16TUfBKwAnzJxth++AQz5v4jtmxErE8BuNdkOkus42n81i4RG
Y5wInjQbQ1nfMFb4lkPpm22HEoMBcZ9DVz4OVzIpQ3NsEpCsMCRGmWcoDma15sJ4hWB+C4fERqtM
kWOGtz6L270jiZksFB7DVtPK/I0E4R2nihvvkiaOa/erTGIIqGQKrbnYXjpX7c3ndOhSJ+SPsZaB
RoM6dvz8n/YBg49lqQPNhUOzKk7dDuBMToKqj5vy6r/28PCYIzQiZJ0fqjf67rrh5/FJzbLxQPkW
6imzuYMB8jGyBFMMI/9X+7Yx0GvmRLP5IOb90xz5zUJ3d8ehv/HEg1EgVCIM0OkI6nn+0D8UxUoU
HFLIO0JLkTb+Jg+20xSigxwEwMvbCJ+1zLDk8Xl39FZCn2Ch3fQ2K7WbZMJkK28zjv+jScCO9DBQ
k5PHUzoI+Hh9Leb8LJFyEJirXoT8mp5BES98wsFSshgc2u7KSpueoloe2MuBpVrOhApMPOg/Z4q1
E+hIqTqhWMm74YbAr8+ytKJ6I2w4KcY6vnX+VRnBdJvQyAufaCFLABcTYxzy93DzxzZkROk0xWa8
QZxpsu5iyWdYv9Xyh07ftvzYte1xdFEC3kdQBbD3j8Qel2fyh8keOzQtPwAmGYhI696ncyUEZocY
17+iLDvxVVyCJTlS8GVRkwHDFzrhgPpK0Ns9c9+SlbhZ2opROU0C/zoCG355V+t27QFK6aoEte0a
NnEnETrkc2Psv0s3DeVFVYPviRpQoX0rMFaUGfX7eKvZWyjIEd1My/83LSj6WiomlTLEbPGhhlSL
vYzML6sEUtrlNTRH3W1Yc/biswn671bT3MnlN03THYDmXxdWOfJ8dEszt+/CsRrWLv0jLn3WaBiC
F63y0d22X9wk5iX0R8ZhqRsrPhuh8sPEcerJ/wgskXDLqSm5pSnP1hLx95WkXzvqZwfMbKXwAOKb
QSfg9EIIqFdQSqKEuTGDQxF6jw49K89nh5dZ0w09eZFFmoftRh+RbKsvz3g2WAlRUqMRYdLhJeNh
Td1fkgvGYbST1s7J6IlycMkiGGG4vWZi3VxEr6j7pL6M0hOUmMFtsQR2SLIXmD4J8D0DGdsivkmZ
twKR9b+LVHZWkg43+orKKBM5rwWNDGBFviFO2rliKp7O4GJI5YyFR9xhbTeuVjyQ6Sc9HJKdvsy9
7tIaDpkY6dQa/hOvh7sKb9TvX11vzjYqlFYqkNVF7q3oXvE7oLF7FNbDQZ0TpmeX8I5CgB4P9q1T
exL34M22N9OYd0+9Z3S3JZg/yBw48QwZEr+cGLeH5dM6o0AIEDTJU7qrigKGtYOsLOZkMy7KUI6P
PXH6ChcTDUPmFMKATHBbnrS0rlbq8F3lWrDy69y8vXvY06nTdaG5MRxxQkvo91f0CJ2Owqyfr7g2
Gsu6irVgEHAo1sM/l8+Hlwi/ahmYumwHctBPD5goLbJah3/LvbgTsNl191ZFnmXVV5LWiqL4x9LE
ExVLFy9GK8dRFz40lFB9LbB7HxvOO7cPAUA5g87LQEIg3gMKq82HH4Cw+R4vpeAbJBUtsMz7bfea
5t4YOErSlmywuoIOnVEmM8znn67BAeJhPAe2WV3N+hYkp6Bexj90ZmNs4qZYAMu6ivUE7/56XJ4h
oxZLRiC+MwL/AgW+1umHf7LE3ELVvEcqlInzDcRW0EMSxMF/wn5FQiI1BUAnqnRYQBydERPbffUq
n0qksZcaXzXClvQfi1rZV3IrXrCUykTLLKz83Xf5y3scEr5j6D9miR5xpjX0fDSks1ZSX5U2wcwV
E9OaaCBiZepc9EB7gcgjKvFMGuOeTNmYYG15XGxKwqU1X5gj80QfMCBSZSvWC5hTkpPyxOVpA2Xm
D6RAeg24hisxG9AqolZ3zwdmDL0fpdeFaBXYYSOvIF36RBk7zkq8nSeegNmZe9y4N1EmSoarF27L
5YgLwfOloztiN/DvZsNNYi3VKfcDQ8BoPm+jJzK4KU5iSg5DSpWcwO6DLgHogFzff63l4/LThmxp
2VXv6a+B6TXmwxIhWb1JIpeL5yj9MWpvol4JwSQlTFKDZfu+VE3GiekLdQ+STSx5ErTgxSO1zeJm
ZmdqgLGa/8lBGoKaqSHptZ3MttpTx35XyS2F9wheBnnmpqcY/2DQAsc7jpjdrITfxfDq+esyj32V
bGYJ4d1Xi+1Fj4oY0ruEYy9B4z1i95pRtT9tfr8LAzrMqFKGYlsIyCx8GinXlsEFTWyXNqrfbhGR
IEXmeUdrXpELhfefaKW08AcMKhhiCKg/cyashjmE3XXHfbF9oyiDWvJiyAMHHd6H4wJrCCz+8QEQ
iJY/BZJT5UAMXN0uW82ZLXym+qTjHL73UliO4xY+YptgMznDDHoN/M7lxLb3AYmukupTy9gGd3tE
K8DjQJO2XEalaOSP4zJS+kEAG84awQ6Q1UhmjQeRcO/oPYH/WJQ64GEbqw5/CoUabrvjLiaX5hWU
KuFSzF3iSNHuqBHbiGSkp/HNHS3lmt4CMgw/Ea2dWFsz2iWCKs5LtYMBzhkUMqZa4m8ZRIAR5kgx
rl7/V4e6PyhLWEM8tbnJD1JJZFembzS3kc7y9G2f/7XmN4NzqGfqGT1oUgIYRKaaSV4+JhwsPlsD
KaXm/B9ACXw72VAlngXNDcUZOW8Sz1eOZBHf9reDzqEbFfAdvYNMOqfAEKwU/Y6b1Hbo9km2m56d
6joyTeexDjzBEKkuq1eISgY677QNHrZuBYI6zClUSvd30ZsoTu9soazUeVo4U22KvorXgn5StXm4
ybNQ7Qujhx65MkR51+WDG7ArkJr/ae5GXm3R7G3Ki7RwKxQD8BNZ17ec1S7mssHJDnJNgfOTOjBy
m+U32BRLKBdx1AwoM+BDsm5WotHvywf1uiksbg9Rka1+Lo3huE6GVHqei5jxzhfY1oU5uTe71Kgz
wL0gnpQFnmNPgiOaLT5B6lqPHoauMdgGZmWsjmK4FaEhhgHcnEl0pphPl05WvDAqtWJn3XUcvONE
ru8JmQQ6rajuSXpUdHECpLt2Fa/2C6Ko+MuuNdYeaC/03HNg6H5lsbW7MOES7Ohq5xiZBN3nVHRE
H7rXtVbJtGN0QecTjLfMm5Kj/5pSA+7g27TJR1Gf2X5BiIk8HlshR+hDUP3xrSQxRHF37/BooiSR
nJ0PN0vLe0J8vynJNc8GXOug+cLGZdeZ2C2ff7sCdKHFDu7RA4WfFQNzq4eOwDDWJK6xOi4+99KA
cQiXYN5EBDifAaj66vqzeGVhJXACt8aiKuo6RFL6Mz2K08jGr3kuK3pvD2RKjpSxMbeC4xZ8MK4G
P4lJk3QxCeFVYbTyJW04XTPG+g99g/tZKSO71zuXeunmm9QomZaT/IynhnsQMUOa67oI/G1oTHKt
4xRofgf5AvGKy4/f+1TmESO1wyZ4LZoi143RAxuI4M5zB076uOInxCmMf2c5gDQUcs2S8pxMkq+f
909CEtRA+QI6Atp0DrH62rRAjbfPtEA1jGBX7o5iN3HbVS2hRN5tpisCteSa2u2XAhqBkAllLgqX
NadqzJSb/jHZKVpYpoieIUIVXBxTKThcOF4SI2tW7e0wNsFxj5DQzQhsIcp78EaPSiAv44z03001
Pm4Pew+H2fGiH5ZG/avE5x7/33pLML6ZVBtPH8uqlSh3Ekyiv9zGWSG4mxDwhfEnuJhjgseIG0Vg
ZDbF3EnSyhzDiLvWI9Q/KwjM5vWjMxhqM0ZG9h1X9JDKJd+giR9vl6JZGTPCgPqq9aQMZbK7+WGW
7j1soVHP6wPR0gyvNOgVYC8lTnrKuZG9ONBao3Ea8EKN6GbcfJk9qJZTGFhi82b1Qj4Fp9Wm57AR
JAquaNRqUFKkO0KzqAqZNOnzRKOQrCbRwdvR6YaCgwSeHeXypZA78+LVhTRhLxnETGNpSV3S818L
5t+PDYYD3XhR8nrxdqBGRHpl9LREPWLsdp3W4ZBdusv/LCAPadOS2hJKeLC0fHtQm0N0ZgZTklVy
wF+o8MJAe3VpKGzHtP4enPfd4xDavEI1wP+g+XLNIPZUO+1u1yWipv+lKI0kvdotP0wx/+A2Nx1d
9e00+dhRE9ZTglr69tTqlP0uvzewnNXFsmQMahncp50vzQPXGfFMxljqCPLlAiQwUZIh6AuVEphZ
9P1KrVkdj9rS2UFxvQa8MGuhhBljAIV8eH6nN5u0570QC8voa86ETwK8GrkXfQIGhKmpmpFIOMgt
UijJ4fDyAdZTcGVpkkk2lXRgMePRfes8mm7W+yLOXXwNXDrModVqF401KRqIyklmH/gOmATVxAYk
0Qsl4Erxh70kPMn2qAmowtbserUjR59EvO2FUg6AYtDULLtmPcaqiRNfumYwCb+2TS7Ec0ewzueM
t4HhZgDHkj2NXUwug5F4QEI0DubdcIgnKI4JByHzI4o1ab/tLRvHJQGiQy0Uu5mALxie0X/t9JWp
pRIfH9YLpJ/zP3kSfHgEsVQqUHugR7lCb8us/pKxq2kiavx56bH28bezJVXFe3jjozNPxJ4V697K
sZpx5xI7wZwfjV63Dn0V1CpXgPR2DbMZ+ZAUvyJ99Zc4OLJLFkcd4uqIRMP5x8WHY8cBdQkZz7ij
Om0ZWqDW2bqzLFJbbs2jnvKf1QcN74fMls/qI7n4/+kr7RoJYBAWZQ0xQv8BR8mwyF2jytV2ChgB
0AjxWryaqVKDFZtKfaSfKWpop3ro4j6XCu3E5KteOGPvQMDYx0btnCkNrFU8kCzD6/XE4XpJTR6S
r9Z8BEtAJ1JI9Grphe0+UQfO9RXoASKTqKsbcwrqnPcyO1Zqe3Sr5NFo1bqj8du856g/eWqdwzhb
7UVc3QZuVFgXcYWn4vxQZdAsk71u5kW3jx5jyirNKnEvcO4j9PNmhzXmJ/W5X7ZhO4n6gvGnykiW
7CmFECkFo5iNGQhRLhNhyGWa8Ubi/9YlgGaj8WVCd1fnI1rt7zsW7pGXxrvtmMzi7X85TY5j3ZOz
I2vCjSZuX7sLuGfz4bwkBSR+gfHQZSZuFzIR++vOQVmmusBGKvmB8uEQ+3+sCX5hnzlQZ/FDXhca
XsfnacvA2UH/3zja6Q18JaAmxj04DTDaVe5YDDw53v46gT/zazZUA+EsdKDLalHiTRPr4lQFXE4b
X/vRwJabj0svQE0M3NCB78f6pfNstU0V8w7DGHypGLPQWXqvXFQd7jMSO4QYz8DOzOToHpJnN2cs
9biEAoL9bHcZmTlIqtePD7tqG6/YA9sxF133kaNug9tz00GkBCpfUgC5PW94jYSzukyQKdD6iDSh
kVXf9/9C1AC9vAPgCNAIARYIf5H4LllKbpW59B7NJ7vm73ZRrqqDIdCETp97mlPc+QyPOSKkN4pX
u1uq5dPUlpyYF1cjW3DEgdifiAK8ymKz3VPuYe2R8B/KAvDo4bHbP72WsXwDIcFqGQarP2XcI0tj
QDIA4MFMecoxSSTdfOXf+Bckx97/Riguyh4pWyjcB8SnwBTCbHnBe2A50f6hn6mHyQs/ZStVU0Wx
tnbycbPuS+lbWQQY9XNdsKMRhD4sbyX7+PUmoepqa49v6inswGQ+QT7ahOVdPFVG/TvG7FMHK/9h
6U7xH1v6l+dSLZGiht0aEbHYbI9msEN1LHIjL7fgLxs8Pa0A9ZMNIM0y1O0j+Ucq7dapjtbiZ/e0
NPehM+oKsbXMcnqmBwkKpymKUj9KaVRasUcx27V++zGfgxtY/QJrWUr5SfQQNhb+HBE2Zv2uve0r
SZ82C2EXS2hjf3PwKsGXVjVqlKMmDOzm/8IxBi8s6FbQX6mf78wWn2iUjgROb+wf4Os0U8f+CaJI
dlHVAXdDce4M3gvehb64ocE1Uc03ynnAr7aiJh0UU1twFdIwiCWFv/ORYhNlSUTPvFqj2sYaH/8C
T/5IRAOJXl088lb0cVgQe3LD+/cJilcHuMpVZGw3uV4veKEWradaZZyYWH8pGZGOp5jWcZZb50UR
HWEKBgHnwk9HpktCx7N8fZ+XWtcHzjQi6A3jdw57rkRC7wtWbzP+GRjSohEJILhVjZa8rj2GPdBK
Rv0LGiYf+UkLjTrTh/kCoVmZtFvrFnxrtmkKBuK/DdU9MKLLyLs3MfXObtzt4I6NBmcvD26o9BRU
hmsKTG5Cchdj9aH7FL2u4gH074IWOYilCCKTPFSvM+wo+JMG2xqUD42vcdF+Mklcia5Qek+zMuUI
ruBn+Ym0eKHefBgB9zciixLrP00ecYtcREe4inp94gWsUFzCxttVLVYFGAR3rRpU5dpiCcvhYGL8
mhZfVw210/x+jxtCLBod5jbzf+UpHZ3C8ekdv8BYeHHmsmT0FLtqSuDSFUbx9HbX8BPaNiB9CkOT
GHIj6w6kLKJyg83IOzYTajA2zBpKjvtCweVdlJ1E5txWW+qXXNyCI1B7+ny+vdC1FkOXAoLmcm/k
A6ESwFtI0HakvY3H+IEW3tFBuFI6ouIJUZExWuturA6fJkmz7Bi++irpKNPCEKmwleC9lwroaPoq
Ky095sKfbmvAipft4x/8iARMfff8el2lOMmIBsJdnO+KKavh9WPUE1UfJzXIV3+uBpttOiHfybgZ
Xe23ICde0K1WHj8RA0gyAr/1zNpQYJt/IB8AMi8w9KSLPVmnUX19rhu4xS5/LnRrB07JD1gghd7g
PbTgJkD73qeSTJbTL/sXc+/QUBU+7yAulgUkj1AeZ9ijfVlSs6tjSxCFNG1H81mXuLIuIeAz9W/e
2Pbiw+DXNiZn+sC6iSCy7Wd3Cmk5Yc74eRHo6h2SEBnwBBxxn8b7xQtTa+N0813AaUl1LuoSnCXm
WmFDvP617F8BgjlGyxMGUJarkeX6IJ87AvmUuEkN+ePGmRgWTVbdCWrfKtcs5RvqBEPhjc1EDAzf
iFsLax4IPBN9DNheSD4vgPuEznDz1DC6qt0MaPnvrWtJqDuyp1e31sxxOJvAGVqqFfBCsZa/Xv4A
QxUiJ1Gh50/7WzRrvKDqvNT0R0osmm/Rg43+NHyo5kc6e+qqzJTE8qSuN/ApDEpgti5cLQD//sHz
esPTNt6vX5+4xZ5h4tXAhRDAUFGIbYzUbOtM43ol1C7KBwAuCIwXvGO0+BqNXIMFMkc1Bjyvwd+A
VyuvPi5ept8/I8JpgicfPVClXOduZ0cXtTQ028xUqp4ZDP1T7cdvsXtDN+ybUZM5H4yzJu6bZvMD
uEUf095tBvPCWMBHWXw70wmgMbZH2eOfj4ztZDeZgsyPo+Jq2xuNwcqnfPEvkv3DqIPZRsNyn/2H
1H00A8UIRo7CRzVCreSoGIS3UigxjnkXpnndhlS8PN5bQCXL/oqgNEXqbXNRfJSwCao6wBAmxR/V
Rw+GCXiWjzcqJrIkpXT/qGNIwHE/0ELCyJrzBlohOZ5NzeX87Di8d6UUY1ulFLqAfoAMbFgf3sbs
0++VoBSH4lMFKwcpC4Qr1cl0y/UukJUzPIl1Jwh5bWi4SMSD3f2Xfs9I1do22PJbKzmrs9GeSEJl
/PQryZG7sXVN/3GQMd/emJXBeWXD30jezBpjK7/Obar9DvXSko6vcugaUSpu14ozIlF+5QhuuA6/
helkoVRwM9El9EtRM8WeE8aSmaZRAhUIw1lig89ysmCb+uii3SCVkkDNQ7iuEDGNAPVsKGFFtqvn
wPbNsB31XHCN2W2AAi4NegHh27LN69yo42R5Xz+gl8mUzTqY6L+Tt2hVZCWQDeT6bXysvHDCJyJO
iayu3o/Cc1IHM6QqAD6MbhPR6FgZE3rKudXMw0XYkyRJ7ydr97+fBLCeTTn/5ijeGD1f8KuQjB9c
ZLfmCGbn66Nd4LF6YPFreadAsbwAUoN5BmE9flKpaj8DCCl251DL5VGxkKYXFf8bJEAIofXI2W6A
jVel1ieLWdPKjpf37tmPHMEhTE6pk6s9OQRlnqPD3XQS999CbMEGSpfNLlU4Tx1tqTW5AgvTXgob
X7UOT5HF6d5PT2FMr5BGWzBK4z+NZTXR55OqyEIikFsmKZN3ADAkNOUXYyi0XyjMKOVYwVRJYWB0
wPioW268ScI1K6Hk9FgDSUUbWobHR0EcOzSOvvoi+vAv77RBoKc/PojX/F5URE0XACZvFtuisTm+
ogN9siFfu/8c7yqX8AqDsG2Msyabl8585lSwKpjxZRIVt1+uOS8ontkggfjpb1PgHkALiu3exV1y
vwZ6OpSpUsW+NW+VTC6S2sozSLwPe9sRH8RZ+swxy6Vvtdpoo0rzRbpu+vXjEEKLCZlBhvvT+MOS
qotEeHjzioLeDD8dwJ90MH7PQ2byXUIKMS6OaP+Ms18JhP08GF0MWT9fiMic635IKfs1pYfgasWz
aiNwWYaVGmDzD7Qa6MbWQWz1FrmYlRQArwHPhy/VWjSPXVN9ytSITbaaD1HzDAMm+9kJLdaukKtU
H2gbaU9XR9a5q/ygNfdg5kYdgXdyU0s8DvUjekm+TSqNshucWGN01T/XpwsdxatKonDJKRAjr0Sl
klRcPTSsqNK6fLt1SQKDXrWoqxO69MPUHfmMEmQ5r0HvKSd9EVF/LYeFO0Kf1L9+KOIAK4kV9s+e
Fj5L9+mKxqu4NXp8Wg1anI4VrhIU4bUZUFGHto11BFo+Eur2tZPAdkMXSeQDesXOVwAzlKGOEYBq
Ffe0SxiY9xTqpRkzd49GxdzkTAbkoQPlX/Zq851fegY6DJdYEVjkVH3DgM520odlB86xnzEtzR+4
5xYvF8mjd4rtiYVu/fmqMH6Nmm9c0X8YIF7mLLLKt4HaBgPr4Fu3q6kK5WNDFsah6CBGzMpfEbkM
Lo/M7OQsNqQktXQamzRJatyTzxMBX2sblQ9sdItZXm32ZPGUU86xc0jqx5f4ghawIWeOOJ9FWg+j
V0zhU9GfmEVOT1hZbHmXcQdBfFbgvwu/AcQ8DvOYa1kSO0UBnXDEIoz4C0PCJ65s2R77swWZQNuI
AjcldP4rU81Bjjza5RqXsbOSoMfFb0G202hmGN84HCo2JwBYOno58mQfwptIjS85kHoRTh/YaU1C
yMMGEjmjmdJIyA6hAwL0OxGqAGvATsNmfcYeYmj871iMu94BWtz12rYVqD3VGs2InjSJozV7uOsK
5qBJ3NLvyNQfi6N3KynGLz/XUsPrkITScNC63877ZfbY3ta/tgNyo8fId62J0IXsAJS0lw/GleIs
38i0zAh00FPGrDcb7R3JYoVnTYV96fEPYXKDW/7xgZ/Qbpi8qfTFz+EZFvjq8yo+wEv1Q2/tLQNq
GU7X6Zfl3yJodaphgiLw8H7dtZxYeodIryNy/KSpapXqTG+oZ5Jri+1DZr+hNZCIlc4vcyKhWF7A
e9mPLWkeFV+UoeyD3tNFw2flwZQhucAXJ8UXindExyaXvZuDTLX+mPPW0NzyLDaPQscChvqCpn4U
jiPifveVm88KoOqbAiqZC24yt8TlSrpTLKmU+f/8sKlPaF7r89J3ISHBpDEcSfOGAPeMiOq6/rsK
3dwt5B5GvcIc3BYr+IvFRSYCq2T+Jx/Oq5HhmeJqfzoQcuuIMAMzEBCpHmo0LCVVaNz4n+xWDFTc
S5ThkJGZE2/HuvdBLHq6TXcSe0w+5ZnFYzzF92uqWQjDBeBjB5hWaA1mB45msFWNHM9vJT8xMjfO
T9IZaK4OWFjuAhDcZWo4BvQFAIuMC49NPUaCR5lAo/ALTeY0UHHPR18YY9p29fX92ydFzUDZu0uI
7KbRpa3B2o7TW71wKUWj6Lrae8IMWGZvkAZDHk6vmj7I8FAo1k5LeAEy/ZOyGlJ6vJKU3Up+vRoq
+TxE90bSVZj7rnDw7bgFgIzxm/iv97AIS9Uz60ZbCD43BIrS+iBQf2nRUCLjuSZPIfaTF0Bp28tm
2DJcmm3mfJIeRcj24m/x3ZyG/3qBOQQHrvL0CG0gCIis3WBUKjZ2tTLfSCYxHg2e4+MPUFdL2/Cw
7dz0fu0tdrB2V7qL8KZ8ysdFqPcUWW74oBqJxznDZ7JN6h+MA+bI6Vry7OUvpwIspUCwIS6qenAR
RwIQg3V1QsoLfZz0OlnuGBa6By4FibggpMmuA7WRqKjHKyLDhvTtKZauGFqfc39DhJzWXJR1bdQk
OVXLYqUIqS7yLlu0gaaUYUDKnZWe+WaOcXBgWAjRKsC5DyO8BrSsDU+oOTYzRQimOjNWiktXc9wR
DUytceySVMbjGqm3ZLPN+2MVHNHTHd3IdGpGo+gw37deuh591vrOnbUaW52yOS+hoGmEDICx9Fdp
KC+7wiYRngk1RCZZk4MwSkbGHcRvU0wiy68AT3llcM4VOEGMlfZsrC7vjzucaZmy0AziEtEE1heL
FcurYuSSjy0RSSoye481/KI6PJumrlk+fCU7Eu4Nsr4Zhzawk5Z80OnyChZDo0D+fNuU4/cngeW3
YYZODH6K5hCpG+ZopQG8fKfZdM8a69001paWfsMVOvmiVY0VOBBcvx5Xl2SwIQJ6q24/C62yqYVk
ttQ1aMO+hkiyzpwx9AnYwsevN/rrRB3IbLQQeVk+d7YAu2MXX0zf7OFYutbVOO9tHWtv4Bqo5M/4
OJdFmy2COAt9UcTa9ZAtXyOXJ4vMXOAUSH4sQhHsoXtpQAeVnU63iA2ETYva73qC77xSE+n+o5hc
FCpcHU+TdsR+KjWfnSdH1m4pDo1nhzU6baV/Wuakj56JrG1gwBHbtWtIIZw1z+B2ssYWfziXAXUx
JQiQa9pIdmlqq+QxNENrNgFHxMvdxfbAe3SybJZbWGLcwxauxDKCT0/RAEj09yHz4BwVq/jf1WGS
v50TVAZ4FlkE4u8PkD7F4KAL/PIn/eUD9o4HUEa+8Z/ANGmXRIckaIrNgxklaedefcLS9UhKhvoE
fueCykJNGJEL944/uzAGFVcWMrtZT/piQ1spd8mAxXx2J3pk1OhIVOY9rxibjw0QELwaQYRCiP6r
73pjYkzHDjWtywmcPmHO0+iJEGKIbuhaBF9dqfbORYW/eZhhT6gUR28g2d/uvN7ueYaT7kZOBJQ2
GcT0LIyA/dmSCCV0iFR94cuoL7vMvlK/LxG3L/zifEHoIf1jah8zzsdw9ppltHm6exmFwOx41YfD
3NVB4n7lmMEO/Z8O5YotYaf+fFB8LWAdXUZQiZmLUL2KH62oaq3iyH56H53aq3IoHhWjMgTQGsYb
/YF9stM6LTpFYIJolj/PpRCpa3KTSFIo5kuUY7I3BWueblJPx8SUZou4WJrrWW3Mq0ruILrEchPc
YDx6J7CtPPv6LkVGRxpTvDPpRH8gVUjmN9AeFF7lQah4P/Wa9SWHmnk42NGedjSEHokeQYdz9khf
e9zQsAZeRYQ9RKwSLZ9UuSAh0mD2xTyAPnxPLNMce8ItEWPksXcNr9cv1RZgRgdj0z5n16qs7XTf
dkWHkFGLJAJCfgqT2+KlcQxe7Cge5vH3bR8hod2aXsaw2eoMP9iiw1mTpQ1ro3BXq4cH1q8fHkrn
C2/2+ezc22CqYi97cth6ThwczA1nHYSFxKZbyL24l1MiszlJdQc7sW9GjpGF5TsvtcDbLctNDnx4
pZZlA/eHQHHkMQ7+yet4XfcES32QJzIaGR0HdzxPPoyHHW+u/ZEiJyZLWR7osnUFqj4BJ5GR87m1
Y+UP54XGtrWIg0g3A4/IiaXDvQYTb8yOXi6W6nm76tmKqpZoJYswkIQ1yYEQVY3v/eH/L1FMiYRh
gLm8bdv1QAgJ27nSgIl9JQhlp6txU/haxxfN7Kk/E6RoEw/LCGGHZm9dQzMRyrKsoWmGwSq3qCos
OQPzJp06MPjafCLoTaPKzZzkZqwR7F4f0oBfU3pTTgl8fjtJasGvwPa/C10R+telUBKyeOgutIZT
Dth/fDtf1u405rsa2mudodBBTGNwGf9Xa3WsEW8VKgYZi8ksQ+7WEXSpjDBoJccoAs+Wq3Il1B5a
iKDZrat8qvt6sp4iE0S2EMNOfFj7sWl7Zrz53vU5nZdj+1L/1zStuB2Ap75qrvw3hFbR85nyK26I
maEdXDSDTd9dsVNeu4dj13oFB57ZXAQ5hng/EUhjzsKOCrqeAjxU5coWxKIBR5aNqkN3Y3Ya1fcB
dFp8Oz0g/dmAg6WboXeGOhHXYbO1YnyqShCSIgktDPlGKnB4eQuyMfw5OXxF4K8rrV7/rjc++Fij
bNXEtnx5UXl+fCdw2nnwkN8kYrcQAqmTFXJ++020z1JjZPir08Fbunmtr97o7qWcVc7FqNPDSywi
0LfPNtAk1AHLO8ZPa4JhimI2dR5tKMOh2IQwla5mxzlcxQG6Pg8VECBdUtR2cWkSsxlxdiw1yJer
/TZQlvMZ4ODThnh+nJiL8+lZnK1K/+zeTqq3lytvwrA+Y5jN605nqnLl1F3kWgB+yadOh4+klrtI
qTQYPGmRbyCdvfc7r+s9Kdv3T1P7ThHSkIItJGWSubfml2TghCACUtKdovZPmLJLAmYQNt/SOLad
fCo7YWF7GTHk35ACuytJ6iXBDHgOhvEIMy+GYTkP5mCOX8zT3eQZ/RDufOOJoXHlbxp79uC5KBsu
tnOMp4FjOOqR2FVfM9lIvvavASsgBtJLqzd4cX+b1o3R//iKE00iN4UceisUmR3Qb4ulgTunXWCY
zAGZj2a+knrZ9mjtUfsf8zwq1So7XJ+Exz7P+8XR5pWRT7l8pYXZGxl+Orh3sDlljA+W2KZSLrVB
cxispOA+0/iF6Nm2CXQFcx/4MWvDmU7mSfbrjxKHszDOyt+fTNgfmSoD6IKGPKkEbqiQda/tfzef
Q92bwpJJtQtlZhfKMRm92YD9ARy+Q6ptPn0WJt4dJZVi2iaYAnRREIdO9032evDEpgf3LZLw6unB
jVv0KwUD+1X9IMKtPFEndC30nkNBIjnH43zAUgPPkU26xfi3o/y7KdBXYQInNGpyDXnqdkVDLZN3
YGt0CQeh4HN9j5i1Ur4W1oLUfG+4pR35Ab/YP2L3KqVLB8s21BkTxhNOHQLf6Tzn+skDEhCvJDfT
vPA95Vz9UIm+80z5LQXc25fbFzZftZgtejfI2sMP7LpwdVGlu3eIuYgqHJSLgmYfyPwYa0KiBXT7
+IXvA/hcM0/ipEf1lErswyx2Tm58tYAgKIuSK5Wd2d+HsxxHXUpabyPegspGI6o+O6zGgo4SH8Yc
j8qm0NgOLHNLXCyl7ETAU/Gi2AaJ7Q6sYGvjCRTUtj96Lf4VY8dc4GosrR9o5VPme/5PwdCeWkCS
4BTgwzdIyqv/FKVT7f0ciXQCjwx8/qW9zVqh6MgvG45yULiOPWhbfMxuFa6zowXcHaiY2CI3NBdY
hNUKLRceKXYtrze+tJywuWVpWJtmDqNTdgnsQMtSTCviovGEkH1bGehkSqq31QkqzKuVg6lwxfEr
9eBvmJ1vF3rymO/oTN6zfQcwgXECiYQ/wpT6EJ0NenUk+RqVGkThxiSVdDcamnHjsLqV8eunTZqT
9h2OyLlVU7k7rYD+u1x0mirhEWkr27y1PKQA7Yq/4bN1uF7FC/U4UZzAoAcSa/Es/wh5JVjkHHbT
i6cWae2XGEZuYU2Fjw3kmDOtUtV0R/r214BAk0KBrOU+pt3lDgvjJb5zfhP7Ymgj/hWLK6Qhtltm
1nicNoOBqPU2ictfFJQF7Pvmxr6NjXXktPZA//mCGUYfPiWfPI3IoZBCKa9kej/qkr4M1wSniel7
jxrOJjBk79/5IHPUqxVoIVRkLL4EFMBYWb71/rj1UIZHbz5TTKOo9KkfU3WT5kBpflbVkwlUj32q
DaH23EuILTEXauuEspkgPX9PxYBZU7eHJs5X0HsiLC2KHYYpreaYkG+kIaXNvapXlKOEJpLOLmEz
TeAQpcwhMCurjN9Ur5v95lrNHXHyy/H2JXBSPhhLJe7MNBpJzje/tmZ6GmfubnZ08jKr/VBhxlXP
ZHlDqUcmAg//ZSd1GDt37ESVz8+igr12QQ8GkEO9y+O/9iydVOLs34qdnhb9KZUoZ0+Gqn/4VIt7
lyC1AmvYFNzfG6UVenTewMWoalqdSDuc5hhcmRpXF0sjLZLPnm67uomuRtjCXIFw7OyVdExvomZy
QFGm2JqyrdpOC6nVhgy4NGnclWjH6ghkRX5gc1xdV77GFfgrfhVifX+1sUzfYZL1RUEmiOk4S7Ea
PmciWk4ehJLa2fFpYXm6kxmCMnVG7BAwkpriFZlUtj/7NEt7P9BL8GViNjoP5DXp4c9wV8WsArNI
XdaqMFQb1A9Vvj8w1nuCvjV2NI2qFFVgL07PsJitzHnc6OwGC1Fm/yBnJZG9dpU/iNbE0UNKLtHR
AWKSeWoAeS07d8gaA6t+HZ7x99Ntg36iZO7mEMg11ynRo+6sfVosyr0R0w8LjI3ejLLQSTjvkFHE
t0/ptT6XKKsdD+nDJQFCU0QyR7PXA6iPSBkmv2GUN9K7ZuKDcza/bTASXlamXTIEMhsMPkGPo9e9
tRi+BqupRADHX5PZFjVYqZQyEwOZdc3vq59fy+12ZPbsUa7R77Ro4/Bxnvkxh96mRz6JDWmRVL9p
AUh2G92EW3S896IaPqe+tAu5QMJ2zVztrXRbq0SBZ6b4mDkMsxzQ42XN7BWI6ncoN05PvDnXSjOQ
+/kJVpKG6pdhWyPPgF9RiFL0kFtaeuFBNK6V5jtKBNabQ76dgD9022JWeI3bQbOOUYHmnKlN70YM
qwLdectQNLauvaKx130kz+266hK+7OJM0OltuIGBMEj2xDqy96v8pMfu4TJ9qnPGVaMkWWkzqj2F
vzL8UbOnhpbRUHdd4zYBBydubDJ8vjFOjk1FZLYLE2TuDVbd6zZUUzWuq2PJ5YPM1Kfc5oFuCrte
0BvGlOI3Hs9P8ARvwcHh4b0+xagoENBbeaZufTqUCNCvTmwtE2h/AA9oTgCxl5cpz1pqubOA26Un
CVuzRbO/Wj41Mns6/7MoC12kYueFc9nd3uxuzm+quyIGaW0jA8rEqYd9QT5hhcNE1PYy01WD0oxt
KJ+r6DqDWFcJGOecLYw3z8aTTyOkV9APJomOkFXwHoHBjXRWdL8DuU/tFJNYqpNTDB/6iwgaAgjk
lZVPzij/DWVRdsdIYOw7H6k4IaHbdHAN5UOhlMPTQCc1HqyRvYiYc93hPm4YzO4IaU/Hwhy09E4C
66vOgNa9gLTHM/HaNVp+btg/EEG48XCjLNohV0TEqqTOdwn8xjseZ+iKTureVAtjiDfNrHSdImf/
gO9Y/LEllXt0yLQ/ezGoWxIeG+Mr++/N2ASPq2oihxzPYaf3kOA+OuyFK4tJCW4nCRIjdrxFcscw
+0T7o/GIiuvILq2ueUOD/U9YbPt4S5s8bzfl4IsCcHFf0lm8gaXI5ycO4AXcW2DDC6XOOklf7/qD
+QspVtmnRFXy6nMI+XKin5IdNbUb8k343nXOCpldWKOWw2S4zGFl2Ip2wRxnKc8+VxZCQMuL4Ujw
FF1ZhSEyLxR75EwXglqv22U3W/IUrcmFUi/TN6BpZDMnghEXZu7gYOEcXjA38P9f3yfeWxv2jhGe
qTWazh74YmwoHDPl/+My50YU99Jo7gp955aj2DG+sZa6Fmnb9oR/WYmZlQLvLUDsN4qiVLZPLtas
9j4nFmyKEmAu+qelbdkFY+iAPf9zhah9XQN0HVYQ4C31oF1gfVh0jLd/89GU8ovw6sNj9IgRb03Z
GOZhSI2raL+65S+DJh3TiEjAj7FIPmkrL2q6KoN4UzTgqtT2YfoMpCefSVr6jp1Oacqx9gziDcgG
O5eNWXfMgcUfZ2oVlSnoIIk2GcXJUKwFDfpVJyPk58u6ivhP9yVDfRSl4kvONXpUAZQOl5tparak
k3RPwMoJOZemhqhhhco6dx1Wq7qK2kG0P5R8pMZuC4S73DYob5Zmi3rMNsHRR9fUYvBBPVjV/5XD
0aiGAPZnzEcY5Cxq7MOtC/2LHWcmFpsjjHV/mGnzhYJ58tGLu8hFxUIIZ42sJYafTQV8pU2Tgu6s
qg8RoHyylZTV5qb3xZBmLjlQgXHwBCPQtdxBLstXpqzpeAISOm4T3ZdKzbc5MWp3gwjfAi9P34wR
hcubS1pQP4FvJHmLjWR5mPsYqRMu6c6GAm/vqbhgB3lvhIZq0mhEGIcRWmHg8pAIred9oy50GuLx
3sLF5MJ/ZZRfz2mh8DXCbfsta1xEb3+u6If3lQ0678ynyAtgg0V6LnFvQvpedAQUsdI9SZQ9Wsh1
z5RF252ZEQomJ6YUG2YQ12qJqElzgrynlT6MPM+F5x7mlOg9QrdCrNZTu6ocK5jSc4g0dQZ9tN69
qMaJ7QJLQie8PfUKvcAkefwiGLq67OdPqzpgkikMBAJGBQQI3GPgoqEsWDyGFc+57Jtd3zFzNqJt
xnKHAW4CS1SK71tY51wFAwZkeuWmqS3hvMLOUIv7XeAA992E5U9NnoW7q69dH6K/F/zyR2RPu65B
KBHxQavVNOYDx/93/tY7WwxDidgnZHHYdk2j4RbdWMt0Nx3DocZLbzNTAptmYYe143quyJ5HJSeg
YGFNkiIh75tog1ILNiumCV5/cNHo/WVVDwRYI4dL36srJrydYMNiMmMk5uctoxvDmc6G1q1aFKCU
g54C9n5fq4nm79uMWiGZrVKS7ULnXa6dL/So4zKKXV+eN0/MeABH6LAXwSBtJC+WLfCOCgi3xl+l
NrcvH1qgTHOhu1oAdQIvMNYDM4XRoK+guW5k5nF2NmxqIeCl80nhEYQkdiMNCpO/YOKABDrPRU+L
MA6IUtEN651emaNggBZw3D76wOrlndFjizPGjZIW8mmEM1tvtagSKXdnQr/eWkbjMh2SLMrdDXI/
P+MIKK9VCLKe2FTBEAyWN0+xI3eAWfm/R+5QEuwMvwd2y2xXuGLrZDFWrqyZ1ZmwGCZYK5oyxlFt
tOO28wvHWd2GWIOgHLm8adKMPldInIGcnhDu9rysepiAtt1dmAAVF608qrwHkSoOPqbmiEFzRN9i
EhVQ8BxuJhA93L4jw3Wuh/p0VSwyA30=
`protect end_protected
