-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YKuQSah0K2jZyViL6RYiSwG6eAAHAZ/YoN8W/6H4jDv+LqH/8Oq1eCrAKY6QOS/dzB87kHyYS3AO
JPXINkB4x4bnLR1vLAW07/Dqphe67sN41mUI5oPzq8BquSnoLnNcr5FPCaH+d4QTHUziZ0L5Jax7
i2TODtb7PQdHh3pXCczORLcVSFLnyvt1Bjn4mMrcnps8DDzVdFfO5zSHwUFd4x5jJ2yjshrnIIms
j2D+ohqrRbcaQQKV9GTaz/UQpQEQZVxbA7U8KxfFVKDoxnOUPz5GornScGC+pOTLgJi83EDSYwGw
LHog4lQkYPb6QzSf6bI105md8qfMROt0p/3iJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5536)
`protect data_block
nGzBP+z7H7rHUNukxm1cbUy4whUtK7OfCpEPLZEYyHz4h0QsvVl/ny7VHbVL5Ire8ZTpzrXd4rpN
sL00Slw80IFi/p9nOZnlCr173qGlUhOlLPnexjNdsmhmWENk/W5IgKWoWaa5aWndh7E6tm8wCVC+
qa8w9ISvEkJRHKyyphNNEWb+C13ZWpCENiP5Amqwj/yAmpQsCEeQLaGVWGpTa+ThTcAnFBj2dl2G
3dzoEzSSFjZYGL6OBf22L16rZgRiafK47OZPM0lP2KwnpsLzx/DCccyF3wlmdlrQ6JcJ3LcwAuM4
sJp6z6cw6NGuzbDI6I+OWC6wqbvskzUX/u/YN3v0g9HG0TFwGAvFCYfvVa5tz0A41HBe0XqdejEi
a5anihKUiHN7y8WXE33RCH19MqanQGofQePufR0kVj/6QC4Z1EkRGAnYE1mCJzNt9QVmyu+YSxfB
FbVLTq+1wxJnOXNBsh98Neb0bKPCRhl1UCspSrQxGGX/YwV1GsVD5JhKwdOlBw5vsB1BDErYL3Q6
Xcc1+IS5KR+RvNVCDg4GpeFLBo8umV3ujMh8rUu36n2i1p4N0yNwzxsxfnLmvooFHfF80bJXZVqi
YF1+K9Zm2wNwVmOWeG0Eke9Wa/NfFu55Z8Cr0C9xfuN8vMcimNACV5uLUwqakTtgewG4qmSPkNEO
gbE4+o5r5OAollh6eZFhXKyQ3MRMQp1v0Kqs1HsoUS4dNM3yoX7F6TGXywRz3Za4yGwSABjfCu3c
HQsva6eYAHX7+vAS1U5++GPb+Megv2BM4vKDdJjlkIk9qezZqUyWNMZWsnmyBUz1eaooBrUuAUzT
XWZ2dZecitQeGfzowVvLRE18Xall9q8bZ/hJZWqW0w0p2Bo3x4vE6bq7B7Zo3hVTycZOwXzr/C1l
uhmE32JRBHR6PaYTY2tkR8s9UF3HOfuW2z9/K9+1gP17VA8Ohzmmalz42c2A16eCLRBo5oiWBHLA
El+3GfNuKAi5ekQ/RxbYUTlh63Np/8aRhAg/UNX6AsHq/J/H46YYgiSpfBX7hFhK93rqKOnNiNNG
0ivdujPx3Hisvy8gj6PwbUuabOf1apVXO6TMhf69Uj3+FSBKKZHkPKhhhvKsowKWtbdYHRQEYajF
x2yTR6cHoEAAw06MFEmwcp+bpi8mOtAOJHSNgEoLUGimXRzywoRVCz8orWbI9P/xWaMFyg4Cxl4v
7yz29DeRB/Z3pq2tzkoIqWgQxbMoERQh9NlSoNw1lQJXvfQjMK3Rf3b68UthpcrWLok2VD6TQQHy
U/rTPU2iPUK1SomCsX/g+m6+D/7arWAhgU3JV8KQhO7bHcIiXXu1wC1mXVX5+aZffaInjYMkfidp
cU8yohJ2HALat/rb1NrqshiBcH2HTAdcWQ3eRoLp4MZtHFUZNLt8raAEBw7tMGoAC6P+fxkoazNb
vXjU33nHXdwnCB2sVv+ZZ/Kb2P0OePDIQVAq07FbyvWNOP89fJizLDsO5M24knqE+xdoH0SNuT1v
h8Bxw0BmoxREvX9GSgG1Q0+bSYRG84MRmcX5sl+abrUD0Gj/CbpAQujh+V36o7CPJlrg9bPJXADE
7hgfO3w9DoNPQeGD00BdRft0LYhb9BPg2dcvX9EqJswXo+hPB5XxHLvigFAugQg5ldWwJIRhhz7m
n5Gd5kCq+srQ/hX2kHDiOpekroUEzUf5zHj8bA8gZMo7MghyKrK5I5dMdfmuUFWQ2s/7rxAjvNMn
0ULzqa5xGEI4xZiaiBvrQVm48wCn+1VYIpNEJVqigR27/WLfAcYOYCh5ZMfZJh9iXJVxYZPrxXKS
UMxjf1vLYrnz2O6y2QzBIFNKr4k5weMWFgCzoYJmXoCDxMBmraiCtDQhWK0ZVryRzwPPjM+CHllc
gGWu1ztubcY28AGCt3tOSxFvo98i0Y0fIqktuhuGddpCMyGZ05FR3kSTnWRBEKXZvxSWKFpY2Qjs
HbVujnbBgxxSkLo2xCeyBzBEo47pOFIK0bRVz/WtqHUkGSOz//9g/Dqi1hY+I++GJOHUmMGKR0M7
zkK8fHhn7JSgdqm+BpUOpSKHmiJsGi6bp0HFEtsnasc9sSr4RmvUEF+aVE2eqM6kp6EaffgQRXWy
NHoU19sijXsXNrWYdQ0uXRHdxuL6zlb0chbZK0AOXlusr/Gn9gbvwCFSzaMBMcGexsPfZF08mmui
E0axq6/M1I2yCjrSvufP2jpY8kOzSA/y/Qh8WDCFhGAZpTHC/Sg/JKDGiI3bDHziIpWeuq7s76xT
jQJxtbF1wYzoIemBfuJAjAO4HMEa+OKWc1BvnfBvoh9fjWDt+eUMrJrP8BzfGgMZEO9HzZDypW3W
VVHxwWD5UAMS2iZ9Bxnd+8NVcBWPwkboPOdSAyo9ThlqfNelfxxA364+qBX1ct85cxP1xj/z4L1v
3wi04Gs54msBMiT0Pn9hATa+bb2idhxa4G30iIYxha/QgcDzB+z35U3NKaKDOzL9kA79E+7m6WA/
z7Eb9+6YnA50eML+uCS/aoiIovHeeR3V1MYYIJaxXhKfji5wqrSJAcfVCgacZ6DzDiYXsRziz4Wa
Dk4Xxfmy3CGlkr76ojRrKNKSc2hiyLkMFycGudwCWrgY3K1EVcxak6thBeAYLqM+v+nOVineb7C4
gPYBqa0HkcC6MsOG9T0tfkCo1hXPdIt0I6mHow34unKN992I3spqeRGzj5ohWnfJGFX3uZMITova
PmPcKrr7fWBCt3DBFN3pBqEtJNvV93GF6QvPrZ7bTeYzXNMGKDkGEWkhuIG2zL1O5k7yUaAd9ngg
Rmda3MHpa7O95+9u0V98ITBZffnwMFGzyyAf+SG9hkYVy5kU3vbetNftgKFLV5OK5c0Qbzf58RBS
mjVpaeUyrxfcjVrrArsruYn5surpQ/7OzCf8TCsw4ZsQlr54YMVjsoqAEH1pIqTAGhe0BX5HeIWk
GH+BGsf4rHGtc3bQpojnIh4R8+P6YCVrNCQlIEy/X0YlpFagQXKxRFnzMW9fDY5Oys7u+5L/2dIR
vqQBwBaRMqROCchLQg5sIbfEOHOqksA78gHWhdMVUKtzXPPaU9a91nStAvqn1PEN2O6/lXmYn0NG
rPTHNPd0YYccJcF8la0OgkJlaWvn1praxSyS7A4Vbf0sQfoNMdiAc/oAyYAe9MKFAJ0ob/jl7pZ2
scs5LhJLDoeE2lYtexV1xwLGap6E6aPoFGu40KTOqnQPdh90eN5I5moLLM7c9P0C2XJ6hq+4pGtT
kdM1ue05YTJ9Hz3h3GHLHRGmrlt3hF0NjARG21Iq8NROsuQMFaW0rjJAa/1gQPxeGPVJk8ABDU0i
0s2nuJGl4W9K9Q0gH3yI48fQrn4N2BMLqyZ5Kmy3Cwu3Y/6jJkjG3YPEDmFeRoJ968aPhgn+DIGz
AbUu/YUX20HKWQoTuGrlAVKzQl9S0xqD0m31TgP+oxPD2UrPusyXlylaMr+M9eLDSGZ9Mnp+dpOo
6wOxQzrcZiPnrUWhqb5JlH/5vqaYirjTrATUpnc2hpxzJM130Kj6KHwFoqm22OBlIw4Pa9pV0GCT
Oe5aPBDu8vL6YhU65Kq7J3LYP0wUiVj/7nbodBbbmuyaGoTby1Z9FlluTuxfa77Tltq2SxwvjLsT
dTJaBy7PcC2tzFENGXARJv8E9SL4IXsRUQ5GJ8/E5K47nno0yhbxRVZzFLf1QtHCp9hzX/zne3re
5UqT76SzmELZLNWsV6MDYejhuUOn+DSJmMK6FlBxgs5s683JTH2rhVwv7VuS2B/pZhyyOGIwSk7m
+KAapVhWNsTdQTgDWQTKUGKis4RNY10bL6ZK7tjvipfgGduPQkc8Qqb6ElvBpT4i1Txy8lUdBeJG
mYhOJ0yjpxyfc/l4RJTRLk13ievgJ+JNA58e7LzyNE45WysPBlfAweitDU1Bbm0r5j6uDIW0jfH4
zYgfEWL085MBp2cJqtf79kyOS+fF3ie4H108X5IKXr+bFz1LQx6MbCAQqH2vkMo70f+W1sZ+wKtP
Mef5LdqqEq1IFXDlX9jvfaWlVaIMLLg9uCesxEp9VRezXSIzDTWkozRxs+/ah6YSCYlIIsvP4/0E
VuhIByMgRIByiTKHw+qq7J0myfkQGTPWzc8ImBzQwb4VJR8WRbKHIxwkEumrLF0TGwJ2PMz1dVYt
v5l+ZsYp1IqlJuqCsGXo5bebMfjLyS6/PtYzlnwhXXL05g4moxtZBTWr8WgQjJOzTE8pPvAJSYyW
l0KLG0RUJD12cCsmY/cYkS8yQOy59ULT4IBR3y3YZkYwjU3MONxeWDQL93sk3e5WurnUK4LCAqbS
DXzPzwC8ro3Y6ulUW8Q4nDUzs3CWU7zuhsYnGiaB81Zm/V0rkSltd8QS6LPPpo9/uI36Zkrg9a25
9Bnpm7ybxrLA/gkuewKuDKdpWQ5WinFiyx/mVtniwznsmOdqNe+3qZlVXQtwIE30/igSbm/PjzVb
SxH2knbykZqvM1OAKVWKzMZ1MJu+PZGtGjpzGBDfjO+Xf5DnukcUhCMHw1Q+uQTfAFKp+KjiYGCf
Do738DpW1oNPl8cS30TVvT/9kq3BcNy+Yp90qWJ4ikh1YHaiPSFEns2V8zzNWzqly6+SI7t9V4lD
rl9SrW9fN33OWT1gfByy3tgtnkTGFRfqS+0sAU6+xJl+Zwn/wbvUNuMihPskXWBQ4110BTOCK/Vx
GQ5aXxV6XjVcgWNs1zH8hJSx3jB1cNZk6zmgN8e0rQTXrWBVczqesfHZrHu9iR0F3nfexwMFCsOQ
ButqPvLlt9vdn5MZA2cQay/GpkiDqQzjMxa0XQqVTLOet/Z3dMoriq+9l3ePWz/2frlj6RKAqSvJ
opMQ0tpa3TiyxgeBJ2y15WpEYFzitZqebgIPoHo0GlSDf00Kscv8IE11HHsSGhImoAbVNfzQHmmx
DV/u8rQUkMPl3NQIPnO4Of2++vByqXKUmsfoh+BwXLr5UeS847RQBuR/H/YJ2kV3eIsabzfqCr6n
9vU7aYQZqzQgZ69UYN/cXvInJo8huANPnyDVyWKwAD8Jbd9PY6ngVe8CBwXr7KHBHo5gT55aAQzv
sX//3DFgI1THunmnB1o80wCVs4NujjnDqYoUezZ9g9j5Urfd35DaxpWAONvtGUe9ueN6ZvCRKmPC
VRmwAm4CFmQVO0niqFqINWxWvfAUjxBRmY+aYX39KT6Re1ZFHtMWLnWGnNgYov0cH50kZUdgKf5W
mvT7BVRo+Lwe5NFBvUxakVa5TH1OvL8Vu2pHXLWtuKQIIYuMFJWc1xkBxnHmf0z95v3hyBnCPkT5
o6ywAgEyZn61quiaUSjeyEuHqehNQiZWw/3AvuxaIO18AX29FGGJueBssCDm+6IEk91u8bYNqkmQ
qH7Ulvw60dCScyjqWrhRdecFCPFsimfVT0bFXAkMy79Rr5I+oLtgohL8+sihgZLYijpBGCUoOXBq
mRfPpskPqiVuU+aigeKvzMZPvsOYLC2Eh1tXEtdLqpbxdFjYGFhbIumbQVZWTquEz75N48jy2WQQ
0TOvxoHA+HDxrduUfC5KoabG6q0zV6tDbHYcjTwOyTZ9pINzZ8/2HlX+WoxckUyBh/mldegsF8Xw
42tkcu25nJsCGryM87a4VmDuPe4qr1DSDTT6bX+QnBURb88hmolGOkzDic3U+LKwaft77Co4oYNi
9FX2pmZSHpV1s9J4OXfFmTS68LcC7+tOcaqk3vbPgkP+hzevxBdN0hNHEj4jZ0Pweo1NBKfCk1Gp
g2S5TCZQvO/CnquymkBu2WQT4qXv90RvdhCOeD3ZfjwslnR8S2wYDaFZDlTnsyOc/91zcVaXrXTh
oQSGKTYblG9PM6ijOEYTFc1irXEh3RqShyPnJElfmWIXF+5Fznz0q4iPFt6gjTuxxjlV6ds+PIj1
bUY+lAOVfDIrtxJbP9t3lXMT6JVi/qkd2uTfnWtI+tIjsWzCDaUjMEx1wruuoI3BAT2p5qBAsaqC
RdBYx+re4n1tEDdSdYS0CbB/7bQ0AgaOFveDPOLyhYnb+1rOPQ9XwiYBztRPgdV3hAiBW4KaRZYS
9B4hUDIf8fq3YZlyGqGrcA7y55V8JmpEf4DHas0NgHtjOUhAi5SDdXlrgRQ8U+OG311P+y8gb3tR
eUoUXtwUnxAZSZClfD97m+Ia2eG6zfA70rgKPIhGWQ0Airn1AL8IGXHrFaFYKpsltGmddZ1uemyG
07muFIXSzS2UtfKq6h/NneODrpk3JbVkG7R4F06mKkc8O9IkFNF2RyZHTY9f+FnVleVPO7gaVqdL
AknbPjXwKTWKtZhn70zjEwfZBiNuRbN8HIPnnjFCnOXQixY6FW8FVU0R23TcVSrQ/k5Bf4vRHh8e
dNYY6pM7CLJmkO+l1+stXJHY9HjcjcKdTqRTG951+rfAbVECK1PMN+qXUD0Nc5kRI27eso+Kz85I
JKtizrz28E589/BeKl/3gJEjpokZ4CUjn8dliNBHlJk76mg1UlBNhtN6OFY3+XTfH7Qvm1JXn0So
2VmsbR1AkcUy+m6udaRN6CPfNjvZZcna11w0M/XLFzRv5+K/sTCTeBqBymiNHt8/V6dySdfCo7N0
rXUbIDvOoCGV3bJOZ1JyDJ/osq8c7CgliiVjn7TFhYcBa7NqsrSlxl2BgIY4uQh/YUeDxb08IMiI
dqZUdMx9XUYZOsSzVcANVsrRe6zmjhXQCNPIVXO5z87a+ybXISNTTKEY58LILhzSY/8sAuaDe/EU
c+KRfGtCj7jDgZTU7JxBSXUwganNo45WElvLT64S/lQFjQ9tzvdaDB1b1LjEKXuwlkaZ+BEYlbe7
dGSuQF3Ouj4dPYb7HtSLZdc3P6EP8FvmxnyA2MWIVdsdToXKDkhaQ9X0YL9PPgF3m/qijcArY2EM
fSvgEfW+JvCQxB9w2J/uZSzVYA01A21UKeobBAhgUjbWUxurpyAhk0A3jOjJJNJmbXf8sHXmoO/a
HXpJ0moMK3lKkjGqZ4slzaCiFWebXKA/aOPgReYDEf4JOjevo+U3KjLF62LqUZFK+1ZAGgjT+7GD
nPgkt4Uh7T6XXKVE8Q3Mu8AQQvppVwVHY5VeshLk14KxLkQhIBsf0vnEHVHm/6xR3k5IHBMXiW8i
mhYw9XaIGvfAlI2nYBxARhoTWp4sVXg9/37jwkrhZGlXLQg6l9UOWz12wXhnBiq7x7FBJJ05JhwE
IHz13ELtozkUJ0q7b/TrA23RA4M5t/NArMAPWiKnIXBxNcUrsetpBvCGNriAM6U0PA4MAz3gF9gR
P7WVc7w0u8XeUSe6vVy0WIilTHmUkgFeJ/xixvCQRnC5+UU2Zo5UMvUMBvqrbRjvrRKViEDkQ/CC
1dRzXFqdpw==
`protect end_protected
