-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yjP+Fj8G2OUUwE+jkJuAmHTUi0uai2+/3EVGcEXaoQlNXWORP0G57TD1ZMlP7Zs9SdHz+KrQwouW
4tXGwKLzjvwNGNJDoziJ5yHj1CElKLmjiAMQY3RueiO3oTPcY6riM/LZ7ba1ytt/daHTR6ufbF9s
5xY6lAJGUDdzkg27R1jiYZqFcMf/5ZNP0Ltw9SOyDEx3DeJ7Dszq0SRyCmOOj/G9xe3suxrmzvir
luT1MOrGrIHFjKtvyQoKp28DxdDUQXaEUq/X1pDtAk9EGMftTmr7/EUSfUW7Ugsi5RixyeviMErU
w5Yi3WExEw3ovVGFm+ibO2GbFAJS4LLMCxig/w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10976)
`protect data_block
Ex7yW5jri7bOu6PWC/f+hrPFDT4mTwnpmEwLjcqszeOSS0QZJnkkMmKPSrrRJM3OtFsokGYdOve7
WAWuywPVbWQLYE1Ij3Z1BHHuuMAp6sK6bm6h6ZTmftBC6Kd6QQE8/jalNgkevsRM06DI2un9PBGX
6bw0ZZp+tEkjPZbPiWb23rXi7XhLMrHKbCaDz1bFrqNxhetN1GEduTGNm2RD7/kBRjFWtlVOz4aA
0dlp5dwxKO6eaXoAP8NCSTLP2FsKuHbQQMgDssH8zIxXUGlU4j4L3jQbwBSY4BLetjUKowux+O9t
LP1EJBqgDRoWRLpSeJ1c/hYcUFCfEoM/zwKr7jlcJL9LFnA4xtkT2ojRAIFXdjeppKRGXEJ/rE54
kwC+MH2pRqCXLX7chRf1+2kkVQAitRuI8q3tbDm6cDWfgtkXA5VrmOCt+xubVSKjduLn+Z7kMg0k
Dq95VjlH6DT+VFFty2HGasb0gi0UQoEJbfMrFDRhMOCBDMAd3YqjF568dzPRIK+spAPMyO+QXq8R
8EfEs2wkMKuCkDBh4U1+bZG/u1uQhTKbXVugZhTX51RVVN9hZ29Rce2aTclcZEz5wtASzVjYgJ2P
1cYBdCe2YSgVazpFMwO4VxhPlZZeHbjWc+05z5fq6X/60XkobJJp7qh6C/8FtNLE+XT4TGghfwSk
06KFn9sBLoqpQUaxoTzfJYz9wgtQhC7rcMtrirLTkAD2Qj9GU392MwYJaogTwbK9MJfdmeDzwSoB
INuV66w+5LLZjSutZrfCd4GtawgMAfaJFpUGR6GkDYU+ldh1sh5nkibKKmwX9VACDOWOqYK7R9ws
oYGKfjSlid7zVV9+axE21XpLJeLP8ECJ5VIvzWnOcQxn069KQZ0R/PMdPl5+f/WGF7y388dyr9RX
xYrhKQDLMiDNs2nHLAtG9UhwaFM8JVqhGoVr5BgL3DCmgwqGGzAqSTBrRaEjzLT4pGhYtLF48mCp
jgKdbYF2CRw1OsiC/OM/TrEN41eIV5LaC9KGC1+9nHa5i42orQL5++g2FZFCdn9N0OmblVfzvnQH
pNE8dkrW3uhrPupCn1Be/M0avu+serJMArNnh2637IVZcOP8ZQ4pucTsGSYtx5ZgWGXPpyvMs5AD
Gl4aqpjCqI1BG1C5zIO3C8q1SNMCECHkIWrAPCf1ikdx6Eqx+4nJ97RQG/qhnHWAM5nh+6+IgO5f
h3WdXLsO31uifvjMMBhUOJVzA8bFuNqKJrP65U/ajE5wUMqFMH/BQyur7LHrjMUL4SWe9mBXZJmG
EASU5zLX1tispS6w0UFWJzWQI7fTDSrXp4g2cqQ1jQy+krYv7lCcCVq9B8qcnV4mdHKW59ccQjcM
PQQ6puZBwChEVMSMhRdAOQJlEV/fECdj/B2GhFOSNbsOGIfaayZwe3eiRti+ztFaVGkh0uJv8P04
WcqAKkrNgCfPTODd2ePCBFF1chYf/NGTzvK93wP5c5k/6OJmQuknRdw7vKRg8nWq6PLdCHKBjsGZ
WT5ZG3vz4EUc5pIt0ae0TB9nb2+mmY5jH9xufLH+xR/kWS9pdd10RWCnxR4iP7Ez6byVqGuGOyzK
DIDaQ4txIQjaOuNFz/w49GabDSjSJOWUe/E3mtSR9nMg+thBJbbIppyloUaY8PiTwFNmx3qifYJf
tI5l7eTpRF4I7fgLSBQcomD57V9GMwUj0hPlbPKZ3vqnocEdi33ka3cLj7LZxnpfGeTI4t8m1MO8
OijMGhsvBEhcPUjASdqLr3djf+dEonzf50/KWBWnNHnrJxbRy4rnFS6LAFedA0N9/pq4Thg22glw
nn+Y1gRD3kJ7NeqjcirgxpYeZ+zMTpqWO9caz+CUrKP7KjNsKItEaFYjkUh8u/Aqjxs3RALp2DRZ
7B/HT5LHaU+T52K7uqGZdPLvp+hEkuD7PwLAtTHW7gguoxvDsvHUh4YXSN5t0ZHN7IjyOst0V/vK
dfcdZ8Q+DHs95Cl8W3sx9wy/37j2cYa7WDjKUgcE1l3hG5Qf3/Bw5+M5chRK4bRDfQJW/S0fg+FT
cSe7GsHDE+KT1c3rep7YFQnb1Ov54EwMwVpIrc12EbN3aZ66iVOn/MdU7gljp2w738P3sMjB77fD
7V4vQ9bIQZVKUexqRblxU1ubWWA0dOaX0xU7VgCmGUHTy013LCNda9RVOdAW6yJxbCIc8CbBiv/z
GJ4rDHhYphuX8wVVk97aqEyXGhTcEB2Risvltia1qGeKbbil9xsul6doChlreN4PkK3zK9mNWmoA
jY1e47IxmsrwStHj/AS9PI3QYnv3pw2901zuZDXEPR6sb2Sn2kQ8Tm3RrXp9JsOqKmUg/0EZf/Ki
2QCGM7VsOS47wocb05QeYeWEUod/SZ3gilFjokIMsZukAKu7Cexh/w/w+aCOh6ICwXSj1Zkui2A2
jULDEzn01amQHbGtbBfpb9kU/JkpVP0Rq1J58zj0wE5HMFsLGp3//gz1ZE1TmWdXge26Wl9dJF6G
kl6RG1H2Ti06Epx4IllE4UV71PAlkoo1W20dCxlY5atGY6w6I/wwN0vau0fygkEVb76ucG6O0BUl
YLfJhQoPLqHym8BHlmlsaNtd/eyjdQUTLkvGieYHxQHJqQxAhm0TrfwLUG6hhhVxF0pjm/HXGGuo
H8Vhp3QNjQF4p//y35y2U6Vzj4KS8szzBIqt+Xtjeu5LtfiFy80gPet4Cd1DBrloyUAPT1hhszwt
smaJnREM63sG5z4ZIMGgVYXfoyvsLAoGPTB2Z/nqt55YPlf2cjD/YJzblvA1Cwjq9y+7krPQjX41
zh7tVWxEN1hZpxWGJfnHmD1gb8SqA15u4c7b+aaScnViYonHqSNSF8AYtn+QnrHE+beIkegjAoEB
7EAAEmPQL6SLxlLX2FLDON3SRAscA7o8wgWOPELyxyVSu2QHDa5/h9OWReqeVT5zY3WJFgKmoYWy
Lq6opQoPDR43FqjFB/D4jB8yAbL9Wrys1TjMorLYKkEQUvLndac6IPnAPw4cImd5mVxgnucqDZbe
SgIyTn2q7u4aagtHPD3OJw4SvUKTWP8JUa6iAF0pF6w0Ez/sSM/1E5UWlnca7IPjR0cgGYi9L5oY
Qqy6jf0sBCgPoPPqABlBlsJN9ijEmO9g5Zrn7bmQZ6SDN0WCEN/K1w5C4gWDut2EVTsRXD5UjMMI
e1z5P8zOFfgeS29+mqkbQfeFvZpOmjT0uciK9jujBWC7heloLZ/PyEM00y9o6dkz+GyavOsNMMgl
0RQG8UsO6s7+LOTRQ47YKY+lha6BC/76niPc/r9SzqDGXxEncR0o1h0d3D+gNOfMXHwP+KBLzhTR
z/GeRNKMLy6B6KRwq/EoSHuceiEYg4CTBrmVVIw6xiSqQuXtuYrvKdot2Rq6fb1BwndzbyF+kbrp
P7kLt/qLRGXpBL0rAULdiDjAVqf55tM3/Fs9tTRYHNw1pwt0kL0aKDIiilZtlvvm62tsLMip6ajH
nPjfSFNNYQQGqVOP75TJtnIrhbXeYaNpOmseIB+ZUO6VWB9c4AYDfGECrNyJ9FWAcOSP9XX3hxAn
KQ9pszd6f1YQ5vYDMLOPP3poyTbJRdhCkGYQA8ySz0e7ryEFti7FXfjnM2qXt608mzoZMzff8+VS
kDYARuhof8SIuNwS+ubL6YDUSYZ3MqHkU7/H10cPTpZS34GzwfZlqSav+QsqN91RreNYqMN2xEFL
pBG6D/Tlr+iwzP2H4ecaV8D8AARiPn2oUoV2xAKzSgLGTsH5grh/WIc43zS3FklRNdsRybW89iUY
LhA4TfTP612yIN4/FMnXhyd7425iS08R/nJqzCYCgODnd3cCrHi0Xs8Fcb5SqFCNZMtrxdCglM+Y
MPfaVagmMcZp/S+295dYksId6+UJlgQ8K1hjmnvAyIt5A6XB3yUooR71hLcPsIPNylhf/j1fkbz6
Bcs8gPMiOmdoshwcSzSEpkMIzuL25dTH3HDgFiHDc1UaA9vjATyRb65XKYCYXsukMho3eltRJiUa
9KzQIEZeuPlCcO7eIYiQ6R/eqfNlokJuvaH8rCwe0M6a4yIndee6sp8/my0lnpA+DFrBbc98AtZs
RhEGNpdE4j1WfWNaRgNfVv+cQmmJHx6vA8v+mk/jHsUIUQxXUVSwbOqunywbhFaqBYCQMN5yeQS8
fW/HK9ZUJYQ1kJsXW0wWSIsHBqnvhQLcHvnUXkGIklIucKwrJlaxH/MK0EttwZCp2/M4DLcMQFG7
rTuFBuG0TTAxjN2PxssVWA+QuvBz/ereqTv+bnJtVwNbvA27HlrdxWVgcj3qShQfulYqGDZM0xhu
Lfg+tPNiJtkK9qEuTKBYMBQ0dm6WV85Glk+LJMyDg2ZYhHzxvoKY+LbbnTePD778xbA51YQRoL1d
5XcPkhncGKnl6ys0SKMp0k89ZHfPd7bANcmTtYCe1hlfipUfWKP694F3Am2FsINr5UikzHCWnzQQ
5Qzl5mgDH1IekkzzUvDgfZjlWoVX74jCT1CShzwXVYD5QjhYt6HHQatJkCKO8Ybi+j2m/rWn+cnx
BeFqN9PKxFHdL0/qX6frIwsnFrMZzy29pFxMC0jbDz2BOBMFIxrIqOs6JsZwRwlevpaUoL2jNp4m
elb4Gt3jO1WVfIkMPzj6nF5yJ4ybzbed4mIcK+d8+pK2r5NTZEcO/Qq3EBKUB3qB07y7/vOT7csV
TFG/GBcbR1p0qARY0M5T7CRaEqqYtxOdcdQPL3XznGdIL+i1FDcETIj0cEE6xst8XGnFEOAh1Yp4
drSb+9XdqzptStuotjNvHnEv5aLDvjDVRplRuAvWQK6L4ehtyHRg9lU+Kgh1MzPRcPPLlhMrxYHK
1oYLpA+JSVT887Q6GYzx6KtXfi93eGroI3cWvkxcdA5Vdka1cwL9X4mes0SbwktvS6EGkDASLJ6I
11CA85ZeNzKqP5Nkd7yXjA6yKJ+whR/6qX9TCDWOySomxvXjmXCD4kIlj9rTCyRH6ZHO9WevTU26
+jeG1ajxwHP3ilRcIIHdGBzd7L8/c1B6AfRRprmS0aIYdWumq+s1hGPrppAjmNbLLwByTC16o5ky
FKmAWiNfIEVaxXOlhlAfS8T08q7PcF1UvOxCdevP7vP8s6626Sc9D3XbueTPVU7BPneh7IwJaTWF
HNxSGGmpK9zHBNWcmOe5HMyfVvBv95ZHgkGqL1Mupio0nqlwN++Y70DMJbVI/hd1X1WcGyAu8RoR
NNZmGnwYtzNuX15kMnBqHmUv0ZMS4P8mZr6sOaFjJWqUbHOkdl7fbOXK17Wo2Ae+gYk2Wloy1xq2
SSBYyAx4r4Miuu2xqRjr0bveNBI3G2Y7K7skUZ8PtWwHAuF0CDTJP5KxmhOZKEzaH7kePCAdJ39k
w7ijLRIGztyT23K4priOS1hXtywVMQ6LtBdhDbbi9duLoKdri0FKbCQKwYEZ2hxGHMp09jfpoDFc
iGNRKiDyWfI2HhdHQOHXfNHJJo3h/8pQoa27Zf8DkL2QLyAG2j59VEUqzmVTYnaV/9RwB0zLwafx
ZSNWOI0KizbEE540X88hIaca+PoIRYZrsvQax5/q1g6JYG/spGPRC7bXZ5DyHlyC0Q7FB47VPezd
JnTUQtOloO3NWbcWc3VlIDClldMqLT14BTJe9Yb9ygORYy++m/KiSf1NWigfSnOxYPRgq6XRv765
cqzUKJdaV/8ZhVC/DNAiILyBWEPBE9sXfhMRkpXr60bAOzLc0qqgQOO5HFxv9mwkU6ga0u56J2MP
j1PXeX/KePuTT80pPhcUmtIqlfie8Ox9FUFURJbDmv6FFzJGWwVP9lKRA2j63yUXdJRMHqE1KQ8U
zfoEtWBkGFLHGeL9m4Ro1mMVvlY9vt7IVvOtXqgXzpMaUB46NJ6A1aK1UkZDfop9negLlfg3uPWw
b+o0YNvuDlXg2W0w0NY32uY/ThZ7Gf9HiS56ILL4DDGBpLiLiKC9NMcyoXSrUjxs99VBVnqtCYae
BaSCa2FaE3AZHKu+IuWCQ6kMBWxWdCgJQ9YfSqomDjNvGccZcYiqSD0EXT9TFIyBotfUA8uIJwV1
BW98SsQ12PMUp2CAaKdGr1I7uvWqBCHrnUQ0fiTZt3/YDGh9Da7hXNL618uEqhVropHHIrUVOnLF
jBTREJSrPQKwN8BbArZtim+SrPkEq8VBpK4v0bNxtZ9rVW2imbpo8ozFniPdrdnOFxFBsJ7av6hc
47seUP6IRFaB6rEAxS6od9XhKdHEkLnibyn/puRasGZEf9RBY5fPIp1ci0orvo0gFaGIep3hsddK
Dur6NmW7uX4/xShXDsaGDhQVbfBxdNkbsoq2rPTW07KyvpF92odrVtUDz3R6VNxfZdrNUX7hUpjH
HqsL+PKXNc512jOVAIp8fOCkeTqwRQIAxvBr7n+wldEvBFQqyUvLs08tBKHALyIwWNnRsuSG+PO5
T1bKyf0BZT+CDCwjIoTG54BTx3MpzZ/OaDEfmSIK4np9Q1kqDKXEJMoOPpQ9d4JrpSC3Az323NPg
AG5XXRy3IIpUpo0YbvAiEQpWpYQS/fwsHSG3cY7ACAtks72KoNi2ttcNt9E69AF+lRKbMPfZPG8J
4VdSpA2RiAChfSa+tLXKUqZKlYwZ4EEsUflNeAtzpDzW/2v0a7tKeym4ukWkFHCqsgoCGtKMc1Xo
elLEj+/DbP7N93FyRcSNrBSDIyjBlVHJPlFTgn2ZS9QC3Sv/MBExTTOOSVWfaCtcbchHiqZkQFH0
M3zVwha5tRl5IufguVDuuYsuiLE8jWmLSwxPEQuaEG63yTDpFCSGDczfcQ8uE74Pr9zRASsSXNOL
ZnlBunFNNnxHymHReI5ek9fmxD/VDbcj0P2zVH+pEtS9Vd1BRdJZ3nTApVMq+o/8+EJTnvLfCvb4
322hjAxWMZ88jzIDku5oi9NMwCW3L+pSFhqItJ1fwyCVrcjB0tjTAAF++1lX3I8OM4dQF5J1YoF7
P6gX6C4x/MkdML8ULUuGbfL+VYbiNE2g81bHpP1bmpgfiJAn3bIniGlYgXVdz1ESQWA6UcVsj+78
P8B9DtlVzTeEK712aqOWN9IB7HgMDf7Zn8nE+6kUX6hLe/hUnEXGhB5i5kpeE1rMwm/K8+5Lnpb7
S9qSlpFIkIuzrvRzeAOqBg8NpfL63gUFHCJJv/vfI3xE35Xm2XoxsPSSs1fFCrmW7sSMVmy7hZ0J
WJzouFVnaN6LMgFIF1hbWgMQaoUIRrJioRxQzD8yMX3/BIj7jTKO1VuvIxeDVq05Yf37/zbFHI1e
M5MQJ/7YRqH/eY66+1YCsLI3+y+/PJVD+o766JWydtQZUV/SeB3Ci9Z4Vs5SqHCimYAD/A8K/4xf
/N0yUaz+Dp8n683lZWYTfa0X8KJWBF3XIPAFZD3Ex+qFtyoWF75wdXBV2Kdn66cG5O1lXd/Jy0c0
JGISajhrxGISG2ZbaHwOIWf75i6/vlYT6NR55oNlRU9vZOdkm0Jhyyc5/Mjte9+HGsSCo3bbN6bD
WNPzR0Nc16ALgblUqgy12MwJ1Yor286ySi2QnjejbrTXeQWAo56xccz/p5m+4d090uBJwJ3RO9eC
vhH340lRjIx1LVOHExWlX3qR8NqSNRZSJeguj2XlRobf4BLR2p583I471qmapIkMEgsUf5gCgMVy
tgGxxRKB53ENYiciStpxQ/aWkd123MuCgsCwXZ3+Es4IK+o/UFXKoFz7ehXVy24yYVV7EkbIpr4F
jGzOnPCCxRf9lMtRQWlxDIdrNJj/YhmtUGoOXMgb6S88IO3dnsbmQYuHpedaIxYfKbZ/S6Un6FmS
MEe6/eXUWe20hcth4SeXnRQBtRmbcXUuJ16lEm8N55PNyp0lBCownp8p3vI1EXZPodcuM7zMr11x
2LkCFgcBnPuWX72oYe+FAkSmviSu7tHg97TZVVj4LWg1nm/x0szWs8YDQx5oeKGoYVLtf5bbG7S8
3w2xvq7cBZzZiHVs8Q895lvZh6zNy3qxTHoQfAKsEMOiOaIJk1qRT33IF+QrFgFkLHl69UtR6hk2
WtE9mNkB2sEVnrFCArLjvro3Ui0fFE7CRAlg2jXdxOfhNsEjrlznGGI9o5N2hGdJSeMdY4DJVJGK
iOAV+uED3kqANp6S6P9ZtcdyTe0gLTHBgcY8c0akDVPnZQIuFjNYn356lwIySuR2m926YD0kDeix
0hclKShyplnzjr9j5p6GEwY+rV6Jqco7hVt6+Tn/ljPwMNXdgb/Kjp+Gb9HuDrN+J18OiQCeGU80
nAH4Q5pOUraE54YPJWjGVtZ53sVWD+RXw68Y+twOGO2KAMXdeouBPFSUZ//Jo3tKfpmJyxy99Cyc
Zqv/rQ0GItS7qMD2mTTbs8zRkDhGqybZf21VPg/tv1uZTUdrJYQhz467jKw+WCWWQdnyo+QEBiUk
WOe6cfEuv/RmXghd40VsuT/L37rs/wNudeqWx2C8FDX9G+w9dxqrX3c6VkUvicgGWN8RXB01iUNN
FJYsxq00bAyXAjmKGAMeXP3sIvBkQWfGf3fZi1UgPGIfbQyXqSy7ihiTz77q9Jw0mp2NZ2k2uSxB
Cr/kIOimBadNYsnDZgeYFBAxMVw+pjf4kPZvwqchGdU7h3/g3a77h+WIxpP+54QNpDupyzXt3esj
lx5/FhlibsxchOOZoggcHgY+oKTtHc3emOz/O7z0WnIT8TdXrU4ultfAbpBugWFsEMYpAIwp+zdE
ziXGJ/dcAzFze7YOK85HU6trp0upsyLD3Qx2mQsPVnMi4R2VZ3Z3/c7+qYfhJ0aLOHoJ8AMKJZmw
M97LpjTcxt1AhvGOzMG8qQ9OgCwWMKYKPiCV+G/0DPWVbwVYy01hc1orX/HIZvvoTr1o0sR2YAsD
y4jvteH+rm8Grjpk4NrNr0ahPoq65O6EVgPJ00cnwNjFvshXqXRKPM99YUfcj069n0SU6IDbrGCh
CTFqDW3y6tkdFUiYydhj1Z1/xGWGZJyIEmygTk2cYfVIXQ9VWbRqKCFIRuvqmsE/tUKTGvcF+d1t
hYxlIstUKsUOfJnrEjzm5Wzy2863dxrL9D/veDiBj4K9RgWWHNcLVRkSxtO/rjFnaFyhZGKeKxwx
GFNvD8oz5VCiKO+DwgvH12kNDOpmfjCiwncKD0mot3dLLnf0bJL5SEPL/qYygQTQPzq9uX/5bafg
jBacUQMx/VJBPIkckIOqtYCGb13CegW7FsjY77ng1pZG7qBuqyXgEQzMYg7Em7GcpTf5I3WqNtti
PEMBNVRfgRL6V/wp1XMhrdShnScuC2EmtkIv8io/uG/V6E27645FRh0XQe4GnpuNN2JXAsz1qlT2
k/GBVgcLh67+hmuR7QPS1KOh2ZnnyH4xXMXk4IQ/zo4GlGuJKqJl2K69zrIdqnhq+BubHJ4jPyFS
VN8qPCJXkKA3rsIbRB0mWPVypw1rwYfLlv9T13ZMBjiqnYgNL0HC2CMgNf3hvn4y9bTOamvkkPHt
NzH87qCkAIZ83RY72pzGPfoUH018GxdL2/MJbg4z9YhLf2kJ5TbAgmlWETwm/KE7+pDaju2/Ok+B
guz9MWso1dtFoTOfENNw/9W5v6hlEW12gPqt75qBEZDqKhTv16uNjyagutGUuYVaIE3ta2UN3ACW
JCpTe/H7RQipkRidkyxMnqxpoHgeQQnn8dvPakHsAg7q40leWxsmOdcvsgg8ITvuThShxCi5v/ex
8afwEp7UVVyZl/GnbtF5BrMmAy21kRyEIpnNt1+xURk+wc/k71RaKnFkOD2YyI9zYul85iDOW2fQ
fCtvvOUaY8JwkHCTeIDop1vh5pzbHDVJy33zAUp4eTCm2BJaGyoFXWDfCOGSt8JMgx3+/7yXhkOW
vB7pcV+FbI8imE/L+HlthuE5Ii+YHb8fOkIZD3GeM9d+uhNSnqoIwz/QvT9b1JYFNXDYCqMfseEa
XzpBchc0rEkS7G/gtbEkhw7U3Rv5JosWUFHMzzS38EAkQZlV97gmyrjNJmDVKhjG6ASdUAzYY9Ck
5h8SjyUV+cg2inuzt/ou3JAjVhk2qnwVPAw4ys2QLXNXOy/CrxkyvoUpabZgBe6LcT64f31K/6+y
857rCdwqq6Hqr/MMno+2xQ9kDHVF45rYaq74lwGTK4/CW3IOY+3xoLLlWJVVNPWGf5XGzUB5vH2h
lIMYqXo4Sa93h997083UNwajY87co1YV7IdciOgwsrpT6ouBbaecO+XCv4qfDW9ZKIrWoKQqRqs3
ViEVNy0XOy1RMaS61yh7IJmcVIRqd6zunklBRTdvpso3xKOMUJtaZQ4xg/RhuMcPmnNQ2cA0NC9W
bVDLpHo1Q36WZO0qgSB3x/35hWM9cWgaxxqZ/NPEb3rwKqdfuraq8sfufFUWX+sITMly9PKHW4Sd
Pk0BpE0AvKHvjSdSRsnjFAgtAcj3H0e0yFYmrY37jT/eXwSdpIPNLC0Op8kua3oXHIr3i7cMGbeL
7E9ydS6k3BZI3sj0GKlNbhHXaJmWeEz/m7pp0C1gXmm21z1h6Z0Ukk5aH97/EAjxju+5VUSIzfhd
QC4KxQBY3prG/NHriZsSNcpBETcVRn7vFcNw6ATBoT0P4RVO4uCEmhFUHgA6/6DwuwK4dgTCnYur
PWB46HZBsq3bOwPqXu99rgtE3Lt2AoGjdBvzTk9NvgtZ5G2msKJpcjDplW977TWBp85JXGo1EEfi
uDOri5M8mB+hJ87uDVzQKdR8OR75PXBbc0Q3h+0apDwbIp7PzJ9LlGkFrOCbpfcOp3yrEhZ6YN2M
Nc980sXF5WwCvDL7Oe+xFrAkJF75NSXFEUGFcJyFb18rXJUj+N+WKrouhXNneNRzU6BJeKQ0AloQ
PZS2vbY+TU0MYYsvgtBtZayJHkLX+1Fss0MEDtiWe6uK90kjJ7IZBeK1PoZxzlZl0wQhCqxxoPPe
vCUUdlvsknCeNHQ9BxEj1KD9T0ihEOiRpc+5JOOqTszSh3hiGddoCChh3jzUzHOxQSMAL7hTlXOW
hU1KU3wbpwpN60wE31/Tw696D5PhlIaTaoAQrKKZFQ9OBf/MeMy/DFxV8PjVwr5+bAg/Ax58HPxf
dw3vQdG5SiDZ/pUet44G7iO2C+/pqyB2J/bYBq4BsCuuS07pps4PNudzME/elYV5KS8bir2PmPKk
5SBfCoRtRuSSTXD8odqfwpa29J52tl+sZ65lVSsSjvzLHJYRLERZMuLL113Bb4oN+YqkZQgLphO0
hnOF+dRwIGLU2RGIk40MjlCh+OtK+yYbzc1p1mqLNxP64o+mZpzGo9G16tEd27TX8zxUcszmHAFU
jAxKkLB41n+gPs8AsrzN8EjFhHInLovDECJOYho6Vstmt0qBQhYuBJtxoupc+dlxoD5QgFGhzixn
FC6RHaOG6SX1dd/f3GXhVeEcsotEHMlTmrIWB3Q1oSGmCXy7vDDqCqT59iHhXz3oiUVUxsjzQ+K0
/HKeqVVUM6fv6ODYig2YHsQag/fsOfM8pVbs9qMFjHaLuuXmm98HogYpSpUcZtVHi6bZuo82plN8
NpjIR3ilAxvQHhCsfUcqKGfolvv0ZJ2sbwn3s1YYy3elefKLSZBxZ6EBeXEExa0z/pMkjddLVXjs
9l1XWyLelQXQUxftpUCgLDOGPC/IbRkHvDOkm20azGyeOzDF9ru57Lpb48W8sIqXqlwAZ13OYTp9
FtcUMF/VvIOLZbZ/CBIAd3tUyAWcvbfh2z9FDyv4QfciVSqxiFxvIGPzRTGHMxEn0lIbu6Jswc/d
/Qsivj+ei0jKVHUdEe7LdgfS/QAZ++LY2hqbReXJwhzdND6wSg52hxx3kKRXa/R03tgtcG04z0EL
zMab56O1UTycmhiK9TGOgM5hnyMbOXWily4VUcbQ2lPAZbk5UCXO0Yrr2LQM88QB8z8bD9dapi83
BN9+K9T9nFnhx/mPK2BOmB6SDIHx+12L8pxGZrrpjY+Q8RLMmh/FMW8+PQgcqks5uxNMHldo7oV2
Q2nDlNh0d8C75p3PfONAUPMxo1qgno096VqINSpfLrjcT+szSf6fACJ60Qt2kisxuE9cnXrfzvzP
CzGUoYdF3lc4y8v6bx9GlYE+8ZCQusgrPlAk0FP9zqpCkFCfwqs6SuBcAK4a15BHpBG0orVf27p0
gPv3y+QqOCLibvwJ/21eRBGL6dAKk7kv5GEc8ikpfgXzRPj/l9jPREEdpgDPzUi+o+dFQ9ZfKw72
z4UsnHCNy3pBXMwOO3jrsrabOp3+whjdcVNTDRuKrTkTWQHcQiVxR3ZBNcfcHprbE5ij7Cp2EXRn
7xQXP8uS2RQs90ylw9hEsiPYQDO+yVhSsFayF/XAXMCZPmH9J/PHiUfO6lnRIAsdpoGzSIz3nAgk
wpqvOFP/N04Zp7B+uqF4sdtHCDplha71b6OH9m1z6gc5waG3BW+SoCJurrHpj4mDSIGw5ToWkJmC
PullFyGkWB/Tnh4rTAZIY8XU+VvT0AV64bwdPBbv3aAGeSwtA0N4UUDge0im0sz798aw3bUURBf6
b8w6Or2ym9ZPDmL0KblG5baKqlKfaiY4H/d9smvwiREKV+TUBjCfW7HQSVPyT0TzT3xsSRy5OWXZ
uInCuRCujWG385u9h6o2RguKza7Tn9aBNsbWhNyg/6c0I1na2LiWBQD4s9hZ0uzDtHMpCj33Fxs8
UFX0V+TFGTGp+DiIPV1fOCU+iVi5TWERiyKh/IN2PEdRzHtVdxZOWFn/14u5OePh6P1uJw64PZLy
qCznaBm+2EhVvgGT7JVY+DlLsMHWiHMHClfnkQNhB/Hmrc659DYOGotulgqEUwL8G9S66M0G+TIY
E41RbNjxAl/ZmAVwuzOUdvaivGoqeQCW5FL5vPRuiMVklfFu3GCxlGl4nnyNP0JF1DqjEwl09N38
ZT/rFzcYCkfLAbc8M+XI6CVvyq9iG96Qr5wt2IM5SgHp6ndSEuK6BqGcmCnLGd1dkRZOrI6BaoiR
hfLWY14ZCnxu0Prb90ANBr3YkOdNbScBMKh7FZu+oto40n9j4lv5ljfT3mRlC/Av66TbrH5xQCZU
JuIwG4Jlybiq1JUfZnaNZbTDVztpJ9jXYwvE2QELC3ChyNxav48d37CnoNHKj6yKN+v67JGoxZeA
PlR9zy6PKUs1dCdxeTDrkj7EX+Z1I6vgPukG6bXxZV9GLFCrvydwzZG1Dm8kF2wxe1BGq/YoHRuf
/tIwnJQhSuq8t1RcVhd1RKM8psQ5uRRRob0/c9VT8F2Yg25DyGZLk8yu3h8Bt2cOQAOcJMJC/oDo
WsIDjp6lo3vSdBGXsIIWwxdah/YJCvUU+QdkA1LjfWNPVUJciwN0Ham679U6fm1VdAFq18kVMWug
yFU/9xAoQ3GgV5a4dSXEmNKyP1j1XS+5YibwxQgfFffks5cbNmnQWXVo8BJdw0EhWNJmQOIZX8bH
FZPvYvjsu+4Bs1NE2vDbwRG48qEM8CDcPuiTM809UYm2TTg6wtWsGs5RAgaz6+gN6Ep8zlLlpO7k
8PpDyyiqYJ4HDgcFDomQ4SWLNEfxMm1kypdOoxjbISd8dimBbiDMRaQsyhAEnSUSpjzrWee8QFRO
kwjTa74LWVl0cdsoaJB7+ULlY8cRp7/2c+mZivHVMillMkgV647B5kXz+1NTJ37089YEeDlKv2yd
98qBSCelSIRmM41O1R6SatZzHhJSwCbD+2nJSP1YY8qxem9aLSKakVKvPPNRhNPOz69tG9iZziIO
ae4PEFoQCFZCALht/FWIG9VShxIxB/wDXKz7WE6RGe3LSIL43tA9cOwU8y4T/wzIcLJNUI7NX9Cc
T7j/+9X6bhXLF7JW3GTCt7K9rPOxb2/58P//YQU7jFgJCZgrM9Eoc0+aPmqbX0Ad3/QVUrhikLxG
MGk1IcmGG6imZfq5TQ5mrqbqfpmsGJSA/DPtSNB1fczKDexPmSE5agaiL8dddafyW5JeN6iemO6r
V4+AlrhuSrySLV/fuAdb4u5J2gj9MY2P/Dz5dkQw6jL2EI11SR4teuqTX9F9e7swNK1goF8yObxE
scpKVDUDCH7o1ZeLIF4+q23imEgncj6gQQmwH1a9nSsUxAW52WQUzywTomZ1UCGTcMm98S8gdWjQ
CCJmgDem79yGRJ13vvvbSZGMC4bQ6UbPzezHGn/UUCGBPQxRJZB0ajLdgV6gp+GALZpN37Ta4R45
dcVMSDO4If6kz9Vf3L4qzWPt5dEn+w+/GggaO78n1f3C6ERGx8pmDqdzYW8u8gIKE3nc5FJQ3DLK
5ANhQcqF36ew3Aelq5udyNNe0Rm1wbO3i4A0GolFur8a6r3CRVwNLBgGErI9Xy3GKzSaIsUzhYNU
H9pJTRd3VIXEiKIQfRd2zPTL/d7HGmnVGRHxcykXvvp5kQhKDSEoEG4U94dKRr8wJez8Wd7t3AcL
xww3QRDp0fdvP+NL9L5w2PX4kIchOF66EizLrrF/OWdD//qH03QqZ2uDRLBuGfrai8LqsZGzzvzv
9ghJUYcgMklwmDKTWGTTfpG+IbQf5j3A52oWL+BUf1SZ/vSpDRRxAk3YRpi9plipeXexiZLs1EOY
vBzjmC0nVN7axolaobMWRFX74Zxi81Xe/2P2a8m8jjM=
`protect end_protected
