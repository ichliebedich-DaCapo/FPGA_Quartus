-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0uXNYBwO73L0xuWoU+z74EcVqX0NwE3ULjqJtO3Hzr0jdiJHnk6yzaT1ptRcmyu6wX5j1hRxuqty
fjfL+Wr+oxgzgCT1C0gdf4RwqKWLPFG7ajiPYhcBlJy7Si2R/SosrhWMb9tuSS7xMKLfp8pF5Db0
AJUYoxQCbigAhp4s+sofMvmSwO9Y/MZ+or4b3/djkav1HiDFqjn9HA7J6cAvSR6skhoZwUUzVx0u
Z4+AilMX6qNICWurGCzM8juopUh6QmyrGeNTczMQo1UH5GMOs+0nuE4UKXMztK76xNIo3UX93fRv
EqHVnA/7gVnCsIXC3f8gK+xtvjxSjNvfkNTTEQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5888)
`protect data_block
kIYZjZTVhxS7M7JeLNxLpw3fwqo05aQOE+18EWE5pmXDN3tWDVvC61aBkcFhyvGgjYDC03soRhd2
uWt2UFujgk6dY3P+3GKTZMN0jrkNgtbpqGaudVLzh1ZIxxX7q5e/DaitFFD8PTVeQulmz4+1oG9I
s8/13nvSD9HXvmUf/oH4BIy/3xQc1rmXic6940nseOdoyIhz/LxX9kx48sYINdlXHSKKnmLxlRzF
HrSGepRYWa4OnXz7PcUUvg/DypLb4FXeHg6PdgOJ3ZQWL3ducKeK7ytvywsUO25qXnu64WBhdhKf
f3rJtCTHbjYBGXvzvbe1rR1Y6l8xn8DvHzRxEXcGSO9RHhE/N51HG8n8++CFURTomWQ/YbDljJ01
OwEbtbJLsJ+PRSQtN7/QxJGv2tsqJGfsARtqJXbw7iUvR8W84d/LmCg3Tfi8yqTMblZZRsHaqbkS
77F+iXeYzrrxFBqIty68xCUOztng1YQNqn55vw7HJ0f8z7o86yaHAHaOzqy8AfDfum9/7PvpvGLl
ATs8Ptq2zMw2S9600uA+9Fol1SK2UWHo0f04AqqAlxpfovNqqlZX/2DpTzZQHzCKzEmt8kHfkQgo
crvpv2PCzTCWRnrQezLj2T+T1ohl7rXnfVvWvMyqaJ/hvOwm6AXTuJb31v4Z5dtAhn0HnmzmRbhn
auSqDMvmEQpicEnD44yKvffQxwFic6H5L2h4bq3jLIDeWcZ9YPw4mfWQ6Te3cDtJEJUzuf9wNlfj
BrdZtbU3JTl692lEa2HbJmj/nYssblZ6HyC+qFXmwH3aJ6mdWCfhsSvADqYCrp6wKc2yPWv77Y9P
XUu0siigKT6XP60zPHEW7KyWQGChc8nVQEaVnw508ErGplY0SCK9PnvhRRdQX9ULUlNtrnnq6m8S
krkhmtMZ+lCEh9myrBoatKNrjxc54nnt+Dy9R9WXc2qwSDYnGMKNuXlHdSGCxMz27QHwoGMzpalf
mrhJg4FnPDh+Ei9R8BV3FYj6UUGfEMhZYeX2gXvlwuds+nyozB19Eb/sZB09Qxk1uOT8oK/dM3aF
hSh4yLKLtP9cgYKNcrSTU5dvJVUVhCfPB5DlKybrJwGazPsCOHz7sT/LJwjIxf6V90OcGIuyHvWl
wTp+8JUPw+gRu9DNXlvFISDLBk3pY8OSfoxoXj+9x+6M1y1D+rr2q8BsTOSLHkeCFxDzUICrPtni
IFK3jEGPxdYOjPzzrBLQT56L8fBqTf6zyzgSK+XxP25MjajWdpW1FpaNS4U33gcCObKdTRC23T7I
V+4tLbEMLdT8Z2E78olnutzXMkzObwGqZP95IjfGtS/zswKCyffBUKIDmszlJWq1vovh9yG9NrRs
FsWVEb8lclTs/SnJxZacyU9IRRnuisfzVYP9CakDdV32QSNLZ2Pj6dF6hT07Fuhzj68zPY5LScnR
c1J+vVOMgo5C+IVEcpl8BLEmEm76PVdZ8IBVDsmR7ws41Ne/9scYXDsjFBV7BirGMM1QEXNYBv0H
e+zryR+SfWHG6Z8NV9JuMPkqFDCY8Yqa3aMd2g4Qxj+jv3IkWPLh9bVh+FXEjIv5zVYupx6oMAJR
ETocBd8/FFYWVxKzyqSLWiclXo1zqthxrKnEt+aSC8SfcAUFdf07/cFJfw/9T4paHvInJ129MYbO
sawqFkIKfEe61L/Eog7+Jk6Sop0cdKC7YU78PHkH46sR3rq8GOW/bSAgaiUt3FzKPnmFpvX1KIwn
kjpr6gOFRqAatjsdDU5MMqTHe1/VWb+4tdMVL8n+7Q+x46/Sj+jskdkQzUZUoCzpRpQZYWM4AtQZ
6QeCTQDbJNq83FzFe3Le4+d06fz+9knTiKKbjUbShz6OHa76F3QR/hkJ3jNKZrwLIMX+Tf37LoKv
lFMGnyGGRuE0PEEou/99S80DIiBX+nU76w3TcFQv9dkrzrfZ2eGhrboFojgQfT8W8Y3IS/VbjPbJ
xtHxX1605XKUXiy6WOcb89YQlXuiWqElzbOjJIoV577F1reUq/b8LvzEof32Q5Ob5ixoqTMpasZm
UMVxdrwcXE4sznz/hSEKJP9/s/8dWROfbAg6eH1D7UIaPgleWoZAHOqD15TWTgv0z3JR7ugkavhZ
GEJ1mWzqwZGjBy/to+QrvrP16dGyPYOH1ud7noOSU13vhMyRYuf74zgh4C+yzOyIOOiOxw+VCtQl
VIuQs5RYLZspQQV5qI8oQL0TMg59Z4qRvKygipOR72YezPVXpRpc9QeivFCE0gGyLMWW9PnOzcMb
LHsnh19NMYyfax9X73PGc7hiLJNZCrTbvSG9NBFAO6xHdG+Ak8x1lMSzccQ3mY4vjnQDtMF3XDfT
HB1L0wJutvy4lc65cA14tSQLNd/x8xcCGdIIMjjgcPIt20TDkhdnBptqpqonDsRIEylzEvNjCQ77
eJeqIhQxulcM0bmDHzdhU/kYR4+XEDLExuvbgrbFVdPBGpSVPQ4/qLfiruZ+cAPLSiyhffBKzE2J
xQj/NwgWlEaB8YZFYIHXwV0WYGFTKtep0GvDya4RMAzGFxNRMtNF+wKac7uA07OAl4C4IpDOHlOO
IqsbhZ33wTb17pz7S+a5pfMm0jl+voKJfumN6kNJW2wUTH57M/pzambAn2yRZ0bb+zrjHmKNr7LA
4owtKmzzJh60NBPfK+6ncrBIJYerEnd8UbJw03N89nLzWbUiKARby3VxTDPD77eXAEYC961FT57T
sAUrG5OHXhDLvDEUd1Zz2CmJkI/w+KdNUNJYrMYoi707800DDglCi7MoGg4jS4rHuYMeCw7ntIIG
0do6S462SmkQAWJl7d4ui41TRWnVtbuWyu3t7s+NirUX0zkBsdNyT7+rTivPgcjFm2TlREjEmLAl
UHYZTSI3pp/Wv+CDnz9p91Rm6+RYkA+nVs3zDJlnPE4CEsleoFGTXcLRPQbjObwN9eMP3cEFazjk
QfFjcP9kKsFja2Gj9vtdisrBy/92AWZA5BwjYYbvcMq1IhQQ57YR65rw8Thzvz/CG9rDHX5luzXs
/1Qvojphjir+82ddUR/eX2mXFac5fOqPSh/ZSX0RnDcS7b/xLU6VpXhQTrIz5GdbBBL9oLEUhhly
JxoK0KEIv0p1NWaZuVSbo3L+scMcoz3u1pTYdYI2/yUNh1/v52q3SuvR+4ZWXXx9u/5IF3dwmG8W
EliABqJpQd4+mMUm8bXeB9sXD97JBsDGAEhUl4oTSdoHiaDAdh1XMwJ73S3mRI4CN836SAE6Q09Z
HT0SyVJui6PoB1jMJSPtXQwbfpv9sG71UzW6BtFUJE+UAAw6jCa/njXOiXfpE5P2bMpdKzTBmFd+
+tfZUMZXo69DwsGX8adMeTtm/giijVrcqwACDccXuAyFqZEU7++FyMZp2BzObhAeteUDbXzaZqYS
9sJb2jTRSO5egqsDAU6J4CYkJZ8rqd4EiZiNfEgKMbx8khh9/HeCO/ejYmWGpWjCRyBQ8K9l9Fnj
J4hyuQol8cogj/QcjhByBt44qS3Ipd/vc6AH+4+fr7rgiSCNzazqADStalLUyGQWKYzHrhmVzwI6
ZjJK4c7vcNgpcnFdnmFa2X1pP/zIqTm0fNho3+p6Qc1rGqkbePbrA+EpiEsPHUR2+0H7jZBNkDSD
OMqcycdxMaBpDX/MmgiE4Uguu9vnHbupoCH+F51O46dN/nfiGuYT76zkWE/9ikjd2ayO92s64ucD
lA1eLK69X54EZ7RlCIWImmFIO6DoJ/NQLABHyEdAH5k1CZL3Y9V+Kr2JSLow8JpuEhk3vobMIb/Q
Df0+s4ioeLmovrRUObbGaAbZnsp1XcU+pd5tsXAhM0ECM6UjQ/jv2PHGiuEtA7zdZjuXel4h5ogw
7nu6uBQT/S52ieX8/MHU9qc953CIwq6c6P6M66MJvZaZMjy3ubTZi/mh//ZvaT8w0KuvmS2S20X8
VgEshH4bqHyjhIOnCqG8r/CMtzVXnJEXYPGjSemLF4sB9bYDGVgfXIzsa3/QI9z51UcS15a/O9sz
RtWymP47V3aNAJirR3mBppv/3olq2tjn99NbAhpKeNng2CSGDyZXkPwJjdQjoYFEx+EE8A6lpo2+
3wRlpM/cgwciEIZOQL9qTOduvUHwqeAJTnkF6DkVQ2SEQwDJq271eWbwWfcXCp8duPW2fdVoiGa4
29z7jyGKpIVft9lpW78mWYtWrXX6+zkgDL2n2SkrX1IKzONY9iL4ccLnH6T2nTVpQ/uD+W+P9XnP
tIxjJ/YyVX3UPbFFakoYgt5J1paQfEqQhGRdGeIA7BB58VzyYvfRODyEtRVQFnuOuiJTBNe+fpD3
w1s/NZ6iPuhiWMlS1NRABnlNVuY2wkz2cO5H1DDWUdJfpadRdeuIo/fak3yTSYhaKPProNyCE0g3
QEnUFasKXNomkn2eifk0zoQU35sCzSZeUV601yhy3EHXfvXjDgMfPcgJKkDQvYpELAR6S6T6v1Kd
5AarZgiZo9PRhki6zskZoJpT61dfWdDE9lBxeJuS5J1tBZz6Dhjx8alfqa4sYBJHklCtenGeyDuP
15adOULKO2Bojq/JuVsRXuvwHZSoRQoYr5cS35Boq2tt695wsATCV5feLWFXF+FKMYZM8bHFt0Fq
KDbJ7m+3+/kj9AeONjl4/PKs+vwIGEhgcKXceuvbQGFLlSoENIlgwdktAe4rI2cLYEydjSnIWB5s
H/MdNOxLkH8bdJ4e4yhNIpmgLBryYZFiS7CyZKkyLuA77//R6wqvJn6adeFBNyhmWx1I8EfziEIG
vHTE+xhET4gL08NeJ7Op2eSCZ/5EIQQqgU2IIinH1ZI4TbGISuyo5eIlcMAQcZZtF+HHakagJmmm
dfboSakce57ETSLeMngLd4sFoWS0iO992A81UNeUEkgCLo9iCwMuxQFOqPWS5QvHhasT84zGCZWr
YSnO/FlE9V836W9pBqOM3cVSJsnHEMwSNfQF7HbKj+1je+VTfBlsrAj8ajAtuqKHuP2Bng0C86t/
p/j3KQC34eC1zk8i/Mkme/2OQfE9Ivy+RHMwe1N0D0f5aU+nrwmiARSFx6icd/GuUvVCMEtLqsAr
6r/vFZaT/j3yG9lrIYjtncdbT2HWujgZ3KaEOab4hZWAbf4PrQc0jZ9IYsgPnvEI6bHSnuV+ZEYa
ciK8TrmrRaVs+rMYJr0XXop6bL7lVCvZ8xnNAuqIo1xBtRIVxMU2QHtf1rKQX09AtmOazj+k0PJB
g7O9zocT37i+V/nPgQFePlFaHt2OzJ50LWSvEW5QwSH+ge/MzvymQaYaL6lrJfCnIDYVzG6NFxf7
LVSnv3OO94mn1JwS8XPTFXXsQ5LqO4EJU2memfm7iErye/L64dv1ydzJ9U6V/NkS73dr5ZbPe2rF
D8iLSRAz4P6aIh8RHHX1JIiKdI8V1JvEhJ6ZoetdEyV5MBA9d1Tu4L9AZck9isP6AODeHWpUA9rj
XxZ2lxd8XoAUmRLqPr4UwGh8dqUcmbfZAiiZzTqMgo9/mEH24+jQhicDbZXLNDhk+D1QC0Dhxp5u
RPc8qKlqq7zj/OLji96rW57is6vJEjaN+s8KCgtyCUV8/nIuCfxPcr9LdFOYtV8TtJEEycnqsIHu
Op32kK1uT+IUM6zB5sVDg7LhCc6gxF84szpYp1uhbTIhji4KcGiBVFmx+YX1H/1LmIa0ICxEDA4q
ry2oQGivi4lu+TDYtEBbQLS1PdayVKmP3WNValHtnaVgXET21/fhM9FIMhUo4pVOWBKu7BjENWj1
TkK0LfcZhHvPIFmhaCafu//X3Qlun4L8bcC1iQ6yb6a9h0qhH1cX3JXNWesdNtodiOEVLJaV8QMD
MfiObgbZtNpylkZzGEn2gTDF0uKElrAemBgd3R6LdTx7q5B/8C3rTTIMv8ML40xhYWotfaFJLZe3
z6YzmaD/BLf0RIX866tmuWHXwfQ3wI29LxgTjdqRb8pWBP4g3aiQCi0xPZ3mcjhEYfxpkeJ4RyYL
gIJKqaj5ZV31QbTn8CR7w/YjLhp5gM9kw7uCcfgfdLHW/82cDPmJRJ99ddzCs9Du4sB2vn82454X
74KgqVDf73vM5tDOK/5nwuDnA8RxsjuSEK7BrM7KdtZ+VwvLym/GsLM7wkPEghJILEnOQCA+IUN7
BL7IT4wcu21XbeaPGHTUOk1JvJHnNC+Alzrj6a5L2/iWOfTagxi9zxRPYFs6mJDWOJ3vwXnO21j0
we2FVmiaYgl/kZwrn+9lVjdfBIudpdbhaqtiJLia5Ix/xumqncNGdF5EC35yq707PNYCTIsCoKba
zj9oAPs+1wwT3ZyJtFz+/v+i9it49hWF7tTlsLpwghVZgJ10VBuCoASJNMhHz0vA2rj8zD2dO+vN
EVIlneOUHuaH8SNRkzOR6h881nYZikUJwvfY3zs3h/qBFE3f7lSMYURlkLo9YgZRfWDLgTpZp6bc
4CH8vUEEIMhVH8gkGZv3mZPx2DkSvmDjv1za0MRWnz4IfCysc7vqCkZ1BjCRp1svd21HchO6DYp2
dCUCrWL8iUbIC+qVhT78mXrSDv+gAYb9gqZ3GF8jPcYmUKYUayeM155uTLfw+1cjefc5RV2g7zP3
3mB/vIKGhXqT6IouFI36n0gsUWOOG+D9D0DJbIoqHT3auo/sfK4l6/dyLffXLq5k0UiKKQebBK8l
+1/cWrnCUpLxn6vcRTUpseOSjMwl4zs0SX0SOCIJfp2UUQpQVfxjrYVcXoBpcUakah4H65rLw2KO
k/UiX8zh3PD2EggiR1IB7PPaHYRSTucu7csU1BC3ohLV9QPeMU6v3atBrREdGRrb/JwDZLoIrxg6
ae3eHn0HjIHhA0aZZUnkew2/iu6qzh62wcBKc1F9LJoEi9FrshLSpiINt5DAcQdXwhaIeG6Uv8vS
8Cv9d0Dud/6Tuv8IF9uGtdShHC9/8MiFBCJ27PfFdO1RYPYLpg8eqw5AmuaGSRG06KMQGkeattMQ
gpfydqRm3vHb1+oHqePz+2q4GMKuxHriXBwHZIhfZjBV//LSevc87tQUxwI3F8cDRWZTMzzpOFpw
9t3ItrsLHL79mX6gn+839ay6/u+nXwil57BRi+eVgijef3d3i3fftgwLpGH2J1I8+YyCWIDs+Ibz
65wVWMAjPjzGLn3DIEqVk2o2/xFY2OWs6jgxQJ6LCy5Bf+SMkYtmCHrCP8CXDNzQcI9nx3OuBZQM
az1nD5MHRVUfvL1UAsxl3IrcZyGfKJKAI/qVuHAB3NS8SuqgbG0xkUqCCqoVEakm61jXEuMZMHbn
JUhiAZbgynwLCzlcKNihF+RUZBsJVGTN1vPSv33TMTh7N6bZTPC01gHcquayww1GlERq7/ut4lN1
J1YGSZT5/CikBcjQizwYMHCkvTQ9ot2ftV9fmvZzNCzPK32Dn7DUYR1jgTZJGhA//UPSsKMbndom
EE+0fNMJuzdjMdHqq2ZcwdE+1v4A5RKlglEQCPQ8gzIeDZchuCsLkVR7Bllz8UO02SCWNpk38EKl
pYKX8PFAx6vCwCv0XnCBGg6G0EkY+oZiqV9x6hIP5wlC4yMJ95s6OKRVqTSUoMjOeEIQAN6p0ziC
Io9GpHuc4UzYftCW4Zy8U4zgPBQOsGO2Mh5n+to8Z5JsaT702BhcNJMGiczjOPuHcLLgm4RBM5fT
3F0hWE5fdLIbYWKCxXsT6PCUbmp25Wxrnw8yxYlpwNaTn0SfFoLsWKwU9CyINj94FVw3BtH4Q26O
whI5VYgWd47NFnIo/ErLMTDPFm1Kd6S4KAmFtz8P5vU5JmUeKhEFDzNXe0h9yiQmJIBEIHXJLKfK
THKW2eudMOJWvUM/xEE+nV0=
`protect end_protected
