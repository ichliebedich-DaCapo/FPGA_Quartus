-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PxUCn2RdPsMKvsflj7e2jr8nND4gdUKMn7ezn6H0Plt+LhOS1ogRQbJCVxpvWq3/AFW9rxMAYPbO
hazF5ejTxZXrDFsjbeNwQQ2L+ld8v4eB9ONOlEQ2fgRBuFcFf3cH4SWmAdt6eA4G7u1fm0PuzenV
JQ5ZPluYCCpG9MB2ji9kSMtrXF7XvWpCFcMm3xsZP/lTwmLApOf4EZnJiW4OBB2fGCBMqYEjlPw5
k7077mSwk+bppTrtHNb9ySgFc7qXlpfzKO/DAtisT4djA7hlF5VfTXITRhkzZHhnJ6XqpSVmDnf8
iwHwg4AjYCBQFB5DTcWBEkW8ArTQMKqP1YMD4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4976)
`protect data_block
L+Xa4EEr6dPQVYrCqnAstnagm0XH+B5rExEmRgXGP17ycBglrl7SsEE6/MPyxjk3vLAv/oPJ7FG3
w2/gKW9Py3nZ7k8P/4mcARsdw9dwBFKDz32aaYxxSkFjR+vDGfGL45ZHd3GDBvGmTnw7rmqlMMo0
sgD8WPtoJgeDcwKFJZrrv9DiUPjaQ0zgvQHn7HBOw9bLwEXiSva9OZgLgjTTaSxYA7S6rEq0ZQ9w
vDAwvWn4G92DLFSKYkdk42EZfAmYUk3Oa3ktZYijdueDHLOCvKJ25upLI51RiqtNL5IGZgfRDNCj
eaKTruSLG+FpE7QHpWTm6UZOl5NCwJ6KuGv8k8DCzMjWMJGb5Fd/fyaSRFxl0K9BfCbzfaO6pon4
+8HdG1t+hRxzTlP6kjy3P5PsMLNAcXyEnt1Bri5wXJQpAE0eO6QdhxkzqYmHRX7YsTD8Qwr4BoMk
CBYK+QEHaVgseaCVgv+oRoQrDMub/oKOEs4jrl4AwdYXZ7evFhVUB+Zzw7tvgDfM8GyqPZ2z5qQ5
JDAls6cZOkJkjNLvbTO3H0nUU0HymtGuzOZakjHF3DjGfWUSejkDjQWw4p5oVlCSWqYcaBow29wb
1BI0K2B1o2gof0nwpRulyjcSPZh7WABpJzSuUGMJXHx4PYCcmYVvmQ97q3poUO0bMuNby91XV+SC
64KfAc1bELclPl9LOG34Wc/301uG/yDrUNtUZVuinQFCZdJfuoH57nQomXmYJQDpWobgcmrvl0gy
J3sZ7BnJql/ITo3GUTuzbk2BVK4GLmDpwpy0PZvERU87+xLj7zB/bj5a/LSi8ObgcmELLOqP1Uad
WyNgkDpWBEyScSbgvEUw6ApqVX5b2mJXJ7TRBn6nBXkSGKRjlGKQZOCW1Uobnf3U/7l1Nb6D9ng4
61FSnia6ki4aw+2kB8/Ij570JksufyGbXMeDuuLzoqz2UJeVvbhsCkjGTkwdxeIejmScVJG0+QS9
tmo31asWKnyY/abmVGW7jFO3d1qD75r0V49XgC8qXJqqVGcODUBd2Bz1/K10a53qHMYtGzlWj5B2
wbuQStRWYuBcc0rxB/R9SDsdpEz9mCqhJorLtuV+vBypgDPoDNXuZyGxh+eNYF8kss1NuTd+Gh9C
227TnYiapQ7Fya7dkRN0noAmh9AJ4oZh25SjPlK+CdaNLdVVZxzR7SeeJReoQBKRDuQAMS10QP/J
U7VGGxFy9nh59brJxq23yKmjOV+SxHP4Z1IIJSnz3p0j+IdgLTIo6KARVqm0Df/RpaqMEX43gMoC
bhKltqHwjg454Bvpkwn4vlxBghfhOGoLeIjwfQuGI8Do17DXtKTWyuL3MFhkssCO6Y3asGuiyxLb
wyNryS8iCYTL+mBt+xC0gUyYh0yE961Cg9Bkp8+Bdg8AV3F5cqS08lnXS3/YL10r3UzpxfSo3GRM
VY16ONU41ssF0tdZ6OcDhHr0843AiSHfeBMoRdOcx5Nb22YgzSSmFH/SRdvEpZ3ohYLbFBjrmdCk
8AkEmkRVYVq1WoKlFh7eWfZ2qtSzd9zHPyYHLNXV7RJqcF6zsN2TPTeZicvXzqwK1iLPBsnk1ncb
Pz8NTrYN5paAfLn6EZO6Mek1pPMhUrN6n/mNW4SpS5dBiQnQGWfsP5iAx3U+XxOmsFMpW0wFwg2h
WLA9yU6nEPJO8zk0YPf9C81Vk1Sy9ieexeFPHcolVya2qwTwuLnerV9CXGVEalcDvelWQ1P3KUhh
YmMKo6Py6fOyjqh6yCJYgw6/l3W34HXHK/VJQv0EpkdKG/bpTlEWMW+ZCEJMlfMmt8FTtR+TIlk2
hkBZMHEVHMUY+bO+3UYs4fKcC/vgwPYr9+SxViY738sazA96lJ8x7UqtxSnihpUF2SKX6oR2QFMK
ghU+6m1pETFqdWouR85RjckSlKwTTrgt7o8SLhm0hSCrjeaxVyRz245EDQBBd6wlATchImJVpNC3
sJPb/RDvkTMIvZNLsDF1C9H1NZ912qDiaUwRjfDThPnljgCmacHbjBmn53zIac9d4+xLDOgx/gbW
2wocixbssdTBCxuNYXzRS+Cy1OHx1EKyzpDP0xYMoOKM6DV1M6vUdFtFRSfUUDBXsB9R9V3EoQUV
B5bvO+bFid55K3Y2FmSJmpCjCRSOtExGBdyzNBU55j3WCR9l/vcc+M3SKOXSmo4HQk95f6BbUKaH
4Jpm/MqrwJIYFug+QxVEg7uSRSs24vBIASJuW2tn94kSv23cOXiVfyVFHl3dQVRofo8rUIVOQL0l
oBBTB5gv800n9oaXoHiim9TYQm5w60ftFYTXn+80nDTmzf8JvTgjJtr0/IqzMLLWav7vtHqrpOjR
cJEGQFT0yI03lhgM0Uvq0YkOX4R7gREyPBz6TbaUqP7uuvaPgEIMd1EGsQfUNhndTm3KIqmNCMm/
DiVTneNblC7lfAcMCgE2VxXN8Oydud/DYm3354DyWTLN+DJYEzEAXldjreMm3TlvFZ5L+iJTvyHN
LHqeyaub2tJJoVCv+llQ32ioY9fURCl9YtryTqPsCR5iNAIVAN+t/3DjPp5/3ywU/SOhGH5aJ6sZ
HHaFNc+Gt8+p6g+eJm51URWVv3BIeywinKSvMrrTMsZhsKrOhQiZnGUD172lFrSZ55IwYSaWm1g/
N7pbicKnm4+Dotvuhg7hOkqARkcLR74sqxEVgEyUbvDOtS5+Ye5dZIktEJe16RYQtxSJsKt4zOfa
X2su8/BL/IWVTX5SWDEmhkzpg6flUzf4izeVpQsbYkY+3gkZirBd3ZUE1HF8hrdpJ5O8X9d+Xh5o
6YC+3d+w0pm0V7019W0rCgLKHVRTMDnLIoGHQZTrNRiwNApxIZKTReZKb+9pP6uzCkLIJGUZCypZ
R08V2sdCJ2J+koWBS7jWhzAPgZZKMOdYVhEnCMX4386YElWS94p2ofeGlcATzVFotoKY/6APx+sc
M4JV47ZW+IXiytW065ESGpUCo95MvLduCN6iR+15r/euPACfB1BqArcDj4kYOLJ5IWPyAaVI2Wvl
IXeKdH6X9gEMFZyOuErjxfv7DhuPJJmiNdFp7mdBhYDkFlCedZUl5h6E4h52cN4bDWTazUoywLeI
+OsiJnRXR1YdbCBDH9N6Sj9hE9oZ9SgypGl7Ueo0owoIpl7KHdJu3EhwCFwqwKmGIyRQoJ6Ggazn
UA2vcxWLoD79mLNeHUgb9sjKd/qoBE7fPIEojFYe3ylkzZFH1IsxcT68K0Q3OUayyYABnCo9oImB
HVCHfQv7V7gUh0GopX50fWPIaYtUmvCirWQbeRyEFJV1Y8U0f7hCpBa27EPErurnY9D4cWyp+OW2
7h1HLnxU5mBgO/U52aXTPc0vCOWLxeKIOsX4U5ObEznVTw4P2Y2YXOjgzIRlGTajjjoQxus3D+Dt
vlM3G0Z99t5cMs7Tv7FRhkCD1GuH8LBEchDJKGwhnCFVnlxyi8sk/u3HpVVxvaPi5nOOcE+FAw1T
2mTflQiGnEhBI0tfqNzet9cV5OA28K1wtWJ124AVuBGfCwYUgYq8c/KeEYrawBNI5JXfmuwYVnC1
Q/xJBGaKmQIOKZ9qrcxfWbTcOvv9bsvgXQU31wv3fy0Z8qlU0Bkf5Jn3Ty8gUcS14sgoKyVBYmZ+
cN17lX++wMLqzxyIkaHro3pww6onkeT97SFmC9x0itU7MT43/IJlJGIUA6bpmHBQCgs2SUtVvzhP
CUP/GFpQNt/RqWPuF5vqt+72TJB40HtTHPhP8LqX/pFfDR7xbVK/mA9tYK+4g1VKfrQs7aPh7V+B
hvyMEk+0JKSNlS70b49wyOC3D5XLNV4vbjyrCmJKjiduLB5NcZZrQJsirymM4sG8DOL8TPRzQH82
ck7xcdDeVW+X5V766Yttne5l0r54JAHhgeHGDd9irj6WWAybPfy9FzeBYALDjtQs2lSKJFtS+YSo
DTaqinLf23Q2ibGVi/3eXNmxItFWTfpFtFW5o6YHtOX9rgeFi+j6y9JyQ0M0fyX+UKnJ7HHq54h+
UkQpXoA+ElWTlIwNSZrfT4kyIhCqnAFKs2ScPJ58rh+SwwJ4GJ+X3Ii4wMiL+9xqnfp5J14YP0MK
NjmF14ibvVv8zjdZlMxxtKW+0y6zHbjOnw0qqTj2NRFi4mw4hr7Shb/4Z84qlulohjWSRZZbTK6r
4I7DztFQg5s9x+SMmY6RdH1vczOZCxsQTX9GcPU15CDfHi5AKpR39jGk1fi1byy7+c481AulJWAq
WvTMNO6i4Yj3jCL1GSdzVypiknUPX3NghfmfR61iFWceBsdQg5JPHM18Au/V8i0Rxs2G7RuxeOl5
jXFGGBCliIl+kUD0Xfx5Sy/XWAvOmvY4qJO0ATozjydMHv6izkwajap+/dztmXXFkDlmlkqozhKl
vpiZdE2evWmR5DfJh7EKEZK6isvf3qvHqfggpJUHVIXGj1UEAZ0sq3Rjx4gQ4nEgRcDAx8Kle3u1
w/+RNNNrmYU9D9hxEWL4dAv0A9xPRKkhUfdvgx4E6NuUOdUMrjx98B/bzaqiwKJ4+1a8ncEP31KY
kI4ECUe4R+MIsZKxKH64clE6neUGh94lOmMmy7YNyw3Ngc9qJMCeJsrKAFKXjU1OgPe4osd9frEF
t9F6rpEE6YFWLGIUTJnNqr5T+LVWRfN/gIEfHFvEBQvo4G3ZZfPlQELcZpdp0VYaTlZU8GlHYyBn
ktn9U63WzrDTncwtuqdb7OLNXoauyFdcwJ3GwX6rf3tMlcJvFp9y/7bSMcntudcZuo2qRUNLxFVN
qe3fssClkFweSZ27Vx0c6AqxaR2obvX+bkxxwrmy8u+WFANmsotOrSC0mKwv32SLnjTT3a3RlXVg
O3g0O/PUDxwfWNvRv0WPSnwlk5MDhKHqzlPITL747AOhs3hGmswAZo/MEzy89m5c1mLtgjxXrl+k
0YXfdsELpaLIekyJYWUDZLelKhos7cO1i/iwMNYGVWQm/hIdceYcxc0gf/n5YW88yJwoTTOad2+S
fVpisSOJMpdefQufTPBLknB6Ck73BSOSSaSls9u6CfRlp/GMFXyZwV4vK8Tu96Mfr0GwD4f55aR3
5CvO/4WhCM9YYuloLqgnLrLactw1DroBM8S39cZdBwuqgGiYBEy6xUZmhSIS3xMl3nUZAw+ecEW6
huczAJo2wAlG8k0sOWbx9KvBOATtGC1JMY/DwtTNaNSuJtXNi8kIJeU6dx59t9n3Ji5SgHPeCpRx
SA5QQKe0uqQgthEoJSl66x2kNmXBnOb3WGcmpkwpHN3O4Q1U0jM+hkJ+nyhnD2WAoEOgRbKeGz+u
apJ7tDQA0hW6+mcKwUqdmEh5GGv/KH9nYbWN0JkokhpdKW6FMg0BqeT1J7YtZfP/xoQoD4iZorbP
QrwfDKOsfHDs8u5RpJIZv1IssoAno5asi2+nxPso3YcV5RMDNSEiBqZ56Tr7lRcExP1KrK9tfu3+
FN5/KRQuI42jhdRf1GbIDk9FQzGrtMC+w+Rt9Zw8FrYrKPUYDRemKVkQGy7RkLkwU824dxSxtrRE
u/5JukfUclAaYUTyDPjAyOsxGI6fNKq7NIh4uG3nL8AwhEj5K+VUK6CXBFMHjnqlpluv2gUckZb9
rpvI63EebBiwi4vr45An7LV1bgjSSGfQxg/h3SVewqt/GazP0zUyUH1NfIeoKK8oxf5+54HO4/qB
uVGu/YrkKQkps677tWfwAvYxLuZfwQaq68i6/z69Ne8KLmO2c2lFj7VIP5YjKKTzLBUSESzwXW8e
LESZqKEOuBiylfTjMrdo8WNLlEcszXcYzhclRGP/RMaDxeCYJ0+/la3C/G/kU6cFp9SX0v0WM935
xazyIuAC0KlTKocSLax86XRuetFYLnaHjOKds97+URQKVE5BdM6nHwV1S1QAdru4ivyfQcO4/LhC
NKEqXU7HMpuL0/52KFcNsN/j/sO4o4HeYXuURf+wBLby1MteCL4atD+u23cEcvtoy84Rl4kLnyNU
dTTdmOvvL1G/+D0Id4aLF5/8mVIt4h8WHghRdFdJJHDIRAqD7I0/uUakI+H/G9cAwATgODmrMyt4
H8S5WnoAaQGq7inxQ9vucdCxJzgV1bozxMnzWmDjckLTK1aB/Y+bYTmgYNgY3fk24yuVyyjw2Z/e
mi6VoC0J09yaDBSgGpW4HxpMyyL1byfjRgcvRM7yOowGIRIlltA1pEmmabjIBGBgT5vIyM0OhgsH
OZJvNdFbAGZes+LCD4oaVM8x5WytKqw/z3i7bS431gRSTeaTe5Md2zbuKRiZQHaNPfWPgLUCTvAC
Tly5U1M2VOYk/yTsaMX7a63qBmV7WFudMDmKgKeKVborjG2YRwwBgPWn87u8tmgCpWGt7s/xFkuY
0MCTchabfqlkuU1r4YaaVn1ZfRRi/k85bBHSmR8TtEiHbRBNnxT5ed2i6Cyc1ax2OSBUxBkRgmXA
bB19+2M40duOCGKrvmx/pbILYjtksWdGqw1UdBLJhenzpUjHJ3exn8ld4PidVuHtjJMwuw6Lnakd
tWT15IMSwYvVHNnemArKaNWLTxSUo8EXypTlYlrkTSIn1S/6LzpuwP6Oh9LCsfuqT4BGwD9W1Gxj
+YY0GHlRso0oQhlt4o/aXSw=
`protect end_protected
