-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZdBwJuEUs/Aohq+flAn9xDEKMZX0S2kNvx7iMaW3HCTjVqFuIPvcltil7QF0a5fEl334sXRThTcG
VYaaOJce+iVO1sOKvAVY9eWs2GUT6Dc0QieWzOeFbEx+HmZ++wcg74AD2N7xv/nuJBEGzmEUNIgc
lxW7C2EH8rUkcmPrfT3r6IHHbhe6xSinTssFHw+SBwJAHIBD6A2FTk6joLn4vlVYDSgKoVj0Z1vG
jguGPAhHnAxSsFpVFDl6o3zy0wn40YihsJsc55A90etGO1JfnUrrLLx4bDox4FcXSvRtN1B+H5kf
u0EimM12dFrCg0htr2qZugNlbSrKvvQENVBlBA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14048)
`protect data_block
pv0nJaMmoiTDsOPh2oDGBCpPcGUFifO8bWOd5aDPZFWcTSBbZAisB4C+8PBoHTe65aVTc+CvVXWX
Ca0ZD+l8AT1YTCW75AtkCrkNDJEmvyJQA/Z9KorQ5WkQGmuHW+5XxhXbdpnxjG8aA5HFq8O9gwac
TldZzhHxq1B2g1aZ4KsV6ysW+fkcRxBFpHFX2JcTtD0eoMU58Rkf+bSKE83RMCqgHjUvYQKRvZUs
QgoFpRiVuQ4vLd3+dKZwsKQ3FxaOVJXjT4X25711RlBZihm9lxZhcQOoud3k+zWiFnnsvsVexdHU
q9FWbsf3J89nAsBYd+1g354zYxizPzWiiLOYDRomQzA/QqLdKd8a7GV8Xu2+s3iYSDOuRuUeSIAe
Be7WkehL2Y1nsqeEqvrr1dTdZx0oiHZP9JRrlcobKb1Gr+AFi/BBAuMR3m8YIpXQ8m2UO8e5dekO
xAYW/BwQI1X0u9XKFYtPM3wpHv++kCdNHhPxg9tXT/AERYcl/BgqmUtBtaSq8CngbaKG9rzpm0Cs
Zf7mAbnVm1XdijAaZKnCq0EBcKQkkuo3ZLxhzbJaXDRGEd0/+2PHZM+e8ZsJ6EAcxxgHgZfifd+n
vTurlSnq4FiJWBZ9n6Ot+zUFMtCoyHOkk56vE4L/lP6VLBQrbgCDKif5oJtq1n/v5bzLXUwXyDKj
Qjrj5VHJyaPDyKSYuPfVCwldN3Ov9JQtMIZrjWjHfFAQnSISoYmmmhHLfl/HbiK98V2L1o2zvdAg
arG/qsQ6G85JGtwQMmDJ6GKDKuAYF6CNLwRr6sUgFrzbjwuAAN2pTPVrkA67LQHVDHf798Ryxt8f
7wYiih2tP2YFF25rD/3WtJGVXIihRuY08/gpqCzA+MRmZ4uWzKY8MMr4rn+T3HPi89s8qIKkwhDE
zuSo75ZlehbliLL9cqvOYtdaJ19ExBSaL4ONP0tC5+2KZbeai9D+YopIBBSuiHT/NteegEX/nSDT
Y6CQa19Cn6M6phQPQPNQD7zajLvVPD/E06LALyQO9LC+XB8qCVt4tfVhkDjH0+icydmBsa345tTi
Ii6e13S/XrytHdA+lVrQxLabPi+avyDjx5JtzQbVY7PaPhITObZ5WH8YNZpdCocsSIRqtIn3JnL9
SEUMe8jxvTOc4s0jJMIu4HdGi5HjvBjwstH1xvc4GM/3udG/aa1yYRmQmT8itUpBqFvu0XVHnkUB
X7L4r7B9s33UMUL4lAuUltzMhW3Y+9mxfybDdpt2YAIm2n7EPgaALhgEwFFfPdNg9QS3Owu7b1Sl
Q2TwXT16G6qpPSNJG/kBJR9MNnCEgdLG4iHrRWI+kLCWckt6bjwwe81QT4HZVSmUU5ze9Wd/TAff
fdY27IRgEQXbfPeyjYA+cvzTnKcNGXAmTwdyjInKUO2h8OSh+rrsfiQXtm7sf58wwfi937dDh42J
Tl3Fma6NSc6yIJHI/h3aI2OcEsOjwvdEXfiBJwJPhF0njvehoOe9LkRrteSW8RXqJbCnEBAUFrIl
RRcKayZqu+ds85jHK7Oh+MIwStcYVbHfVyQzHfqNrf2Dl+TuPS64YnugMPi8O0qGWPkMzrp9FZBy
pXRQ2STYgxCRaazc+HPWrAFQhuW4rT4+pAz+aj3JBcBk8aKsss5osNNuD65GgtmfwLr6Cw4ZU1y7
+jCxnzxZlIyh/Dww99i9AqqJPhtlq3GBnecFjj/abu8l9C4BtO6xHd3zWWKUwMMqLVg4l46AjCoF
dyNW2obyRsRPsA1OiwNbPrCLpxG+GMw11aF/rDHhdfDDM7qzt9MjpOGLWm4TdDg58Zn9kH+94qKv
W1o80PURN+qtoBCZvkwtQNi9I5cZudp4eXKPLi0cQN1ttrZ8TcPrmhcfv3oMSmcX0e07uRjRISr7
0ZpUOxbYKrdV8o7wbgHtXqOi5C5KFEIMs8e+E43cMNQvpNQttrKUST8RAOJUGMyxIqKHK3bDQD6T
HAw5ibwEXGXBo6Ri4Do+yrj+7rMw0YdT/vViwE5mqo3pZMY2n6m/sLw0JK6CqCQDhxtFu3Y8n6ML
RAF24isERYbs6jp230IoZkoUQEoEycrU8Gtoetq9ssnisBy/W3+cyOX+nI9ETy0p033f9dJrcdaK
wNJq8Fsi0fq7PsU0+LmyklJzo5ybgkPXAyDOFV7TO9+iivooFcAFsmt4KEHli4Dchbwb9R83jZ0s
D/7pbCm9QinVi2aSwY5RnXBtKGb0rDArM/BuaB8NuCzQde+ahoYXR56pJPHdQf/9q+2Hx7ruTQSo
0VCoGd+vMMdwDu/avsYUIzrg2dzWad4Wg0/qJIB8cp9mbWYY1E9FEtpusQbO32gRzzT/BKxt8jS2
KrIcnePb165hhsphJyRTFOZv+/Cw1encHTeRV3gavmMRwzkRJCIA1/VvnPhDNM6D5/+bRnNxzmUi
ZqFXesBAGMmZ+s7eQLqK/fiy+ENQZsg1bsiKZNj33uvN+DD5aeDClZm3KJ0/x9q0MxCpennta6iX
/HAS77ff3izhswm0PIEWbjTF+x/Mk42QfsZgd5pInasG2YtWMxtvFESVTdXtZ+nrHVZyrhGMiCPa
+WQCN2qFiNYqCBPWm2jPE8FIzI9UIMGB5zJZmmkwxz7kuFHUayxOIuBy/ujo+yLzyldvGGti/49t
N6YVb6YWgQ5wWhKoKWKGgGQsht2HQAHV8Kk1IUCQb4e18oQaK2qC6jnGYtzd5jUtVSehgbAGdx5m
p7Sva2vHcf3r8K/hHbIxfStJEvKYQWgE6+hkJyrG/CH/Eec4mUxBysamPbiUB6iKpSBldZu1OSiJ
w1lQtSJHbMypuSogCC/WYoXVY1UrIVkoQhNf8vkrpA1Np0tk49vz4dXaUKLgF78GHs9/PJZwuPdg
fC4pRpwQQxoYCmMD/F75P1wzU1gHqnl36gSn8rol6PQHZRNhYPdNP4I+ZifKp1eOZUChEGJLwvD0
Tq6fvtW3LpWcj8W+3LuT7Alz16hWjfAwdB6sXaCDzqHg/d/92dtKTWleNU5ppYG+6FRv7BrD7+qk
QDzk0VkRo787k14ASPI30m3y0tadeiyoPn8ozaBfexCGAv4e6jh9gNY1xS77+aPTxxCVGgxR2IUG
Ep+x49vUu+XiXl31nfEhZXkCMhEjBerDeKomLh8e7+Mnm3NO1mcTgERdZ2C0SVx4ktL9M3F3TdBJ
JFqfPpIrzgnK1njxsB7xfFfgjnvv5tyHdmZm8gCA3rEcogmv0AgWQPm2Q9VALeGs74pqTTvXzFCG
IeK0FAMP3sFilpQkK1K1OgvB9TUIoTVWKT2jEjeOut+6ORGdZtuxJ7AEyCWPkYhmV6E9wfOhJfot
NZO2Y9GPScIdhE1/9crSjKrW3tJs9O47wFu42wA3tIhHQu04PpdfAH1zY//cwJWN3ksgcqHXPCqd
h+Sj0ACYr1Cvnr8E3jXarA3Zv/D7pCpCKZC75FtNmuQw0IAxQJI34D/hJjpxgZPhE8oNiVj5peUd
nycHFG6pmGKjuhHVCBvZBD19gXaj4GqaAolzcShwOlt405PW1keyKlpyOvhMns4OwUfkx6Qzy85d
cgGh1edPHlLCy+8biiMEedgIuf8GRMFIWGR8VhCzX7TqXyMeNgYIUZHO1veoTzZywIYN/pVmxWMq
f3KaseRzS7PLALBxe55K0Zax3L8bTkkst+0niLa8QsJV9yugtYIyKARD4BM02dLzRgxRHGZrC1pB
bnThUDwlrZZQAeNmneu7+Y3evHqpiK1Z9N3wy9y9shkWOB1AjA6fEccWw8W5xLmSfUAXX5Fyxate
vz0u6ZwxkbyFbIGNpAT9QHzxOhOY5M5DUpyWOwahn1TL/NQDCp5uKZP7yG43PxdSYBGfQL4dOZGL
Ycei1MtI295PbIwTbkGKh7WjVwWthoN97Ve/9tjmcBfMbSI8yuQ924EFL8Vy5cQLuQdFaZfcVkGB
iCkMs/rUJangZpCCkhBR2jS+BXafY3bHAUiYfyhhFpSJS39G28vpPzNdo23gVgLc4Q2DtrdYNrcl
Bm9v8xmydBD6qypqHoPXJCK3uQZ+BYIpDoGmb/ZeKVTFxBW+aS1lknUGwogG/e3DpWOtIkzgaACW
twcKtwwmrFLLRC5FCf4C4jYuH2uXFi3qQf232J/gh4sKyJKmhJvh/ziWyAuraU5e9BIw6L0F2xIC
MImqdh3u7U52PyEmKXjabtYHrC7KGts9umn1YAle6JKe42wbaUE5v4k6QZ9siSQWQUE8z5KvNg3q
uvaAu+XuiKqq6uTjYKnvP88QFaY26CsPmJf7ekOfwmtb/tEn+7U5TJXJcE4mdO0yMMz0IwR2Fr+o
+00xx8NRgacX/Zuh8/1Tz1niEzio7fHqDk8N4YLY4RMN1CpnG2L3vDsZjx4G4LrIwz7FvXweOfiC
MmTJCOMf7QVjPhtEnM17vNDx2C1eMjJrq2df8imnurciBzRrCxYXgT4I6B2ilB1kRDD1p1cUX8iY
Ff1r6yN8C/h8y2LbIEOUVXG/DVDn5wAJN3sTQw/EA7uHkR1Kn7p6rkma09fAOa2gFoIhenzNxkF5
xDRdP1eXpxOGWwVjQMORJ6HD7v6mp3ckijQXXPikzEOR/iyn3eI6KDsHCcw65PRMoraiUgCeyf3A
4VW859tKcOuGwI7KGW9ACT1HAiG3VxlAAkzSybrZpXkcQ2xTqroWADnxSh/q82uZEHJZmNkxcPJS
A/+/NSqKjGsphxAOHJSyRzehs7w/RIiYoOhbQRqKoFgTzp+JApQLel+8JJO248u6ggkJzNUadDIx
uww/v193aAFvOfoWzFDCEyQ1Tc9Z5ylE6nl4SPgMGhEWUkrtMNR0ZSTabXc9V3KLI4ZBUy0uaUPh
ZFMpHKkj2DWLT6cFx+LLi5AaVG1ec+/UzbA13vuvXcw3Q3Dvr83qJtk0U0aFTIVVlGXUDYQXH8/g
41Pjz64/LQp7+A7bK3OUcJ+YQWt/2QlfBB3CVwvZY9uPUMxCztf2KvSZFpC3N3EAlPDR5nqLGOe9
6zghRkOSvkj6E8kr1m4QwduNAsTxUYCoQw2V2evAc8ZuMXbK1o9ItPB/x4zG1/25QyOgAJimS7U8
MGinsemaBySZQ2KJUMYuBgjO1dbhDGMrOXhVWjdUKz0wG18eYungEWmMRtI+jZF63AQ6/Eq4JIQ/
Uiu8q2gToj1EV+uZALQDi1m8EYuifvpaH5er5r3BtkgveftKXEH7MLlKAO5PUfK1iBzQgzXI8xLG
vR6aoJIV9x6RBjuSMXd4aVaeQSUh8fKzuHMVV1VWeaBgSHT5sfUKXPASmNn/BGz2ZKRaRRV+Kizt
uPaOM7tV+PoMooquN/soQBVSHjQxRmRlCrij+N08gNttr124E+yYaG9v1KwxXbUZh7uzQCrC3yUY
SnazBh9GlWmvMKhDj35+gNebATc5RYRHyqKHaOMXa3UoMs7qRTc51QnqARw8v3KpJ/WWsXp60gyK
LSOx2o4F9oF1Ail/4fGE9nsnP5FC9hNTXOHHiFQJDoKDIEaX+wIPR5Gzv3o1SOcmHfasr9Psi1eQ
WWBI3tMfb3DLwch63ACOW0gL4N8KXoTIfnHLwVldsTI5fqK1cZF4NU6rTDPKNQU3NZyj30SnRuYD
BVxvyJ7ssXKiuaB2h/jELly7qPcRNxseZ3GsT83r/uuyVwEOJnfpStbrHIbXLY5GCnzEhx7/GJ3V
pjiYkHcq6gVnSXUo5pS75zH8JCrM3IikUcmWtXSjcZWGHiiBvYo9WUHOhMtERabiHXthUje0R4rM
C7gSWvlWM1iAY3GcZGz5kjHQQPCWLeUrEtCM1PEIgCmF87AgAS1v8t5CtSklg5lFBNsnUJ9YkV05
hmJEv9f1DAWeEfSHS9t7IGSG0e+qXE0zXjD9uyatldns8nTh9uiCq9kSO8t7X0/wiFxbEw82QsUh
nwIZUmSUsiq2GFSN9+6V2fOAuoK1TllJgR4baw6cggTlMXNJbFxIzMNAQ6lKryCe/RJbUNlvSaBs
WDKA91u9oDenT3D1XqwmMzkDVuaVlVXetLU94gaSiel0cwLwCFdzozkVqsN7YDNC93Im75C01/yH
v4TOax56fdI0zkx6nbiOIoPqJRw5rmIpvwIBvg9nuTOXt60R0CXzWt66rS5PYAk0glJGEPm7leGG
WnH+8djrF8kMuJoMoLg3U5m8QSJRRyv5EXoQUGF1bXvHfhWTLx6BRFuU7zKt9iNa89eO3FQARlT/
KVTEdIYGmrul3gI9RrBy7goisXy+gzNI9rTCKZKJCbH3mCDoaKzhkl6x/CVDb+AwHkNfHr2LTw8Y
Y5+7wq0Jb5eueE0VMvO7G0k+i+3zJ/zAJyhuC8EBSH/OhJ3Rkv/Ec/omjM7gGdgGfjZ+/xFE2WrS
vsUg6mVY/argSphcAr/+nWIjFWW33O69rdET6w6WprgzmRu7uUYecFsAmAmoS8oLLNehXH+64PJM
SWmU/5ynO19R4cvRZH01ncd6vzw2EEJu+Nn9DIv7HV6h57cGQGUgPL3Ry7GPMTSranBa6pXabFoi
bhtpaHuTuau7TmtRkBgcl7pZ7Ng6q+qu66hmfqC+WY+PxPUcbMDnVx6k/51h1GKH5Ld0UrITj7Ru
0rztTxHI3obzuWwRl2sH5ktZN8FEHd/RsP7HmoYJJXzaG7Wy+kRTixHa2lCW52La8O29yHNMG17N
o3z3Kej0lZD9n85BoooOR7DSRNbU7TBmcIinvx3jHBUvt8R0naMb78UNqFcjUtDwEpbx9tGtpA4h
F5Y15zpp6O/x0SZ+oZqz1LiDmDv2FYpWMj++AAafwl5Sfofxnoe7MLNBBo2ijlvC3pqWbK9Vogfg
uznrJqvjnXC9obVNIldOWzjX89EYwGE9Gp6e8hfCNG2oAOv49+VWL1QtivMPF2bcJinaXtwI4va2
5lLSuI1sTmYCVNZaBT7HPZOT2uv0P+nxjdhH+jbWIvkA3ScNGGLYZeROtXD4ZAE+6MbSI+NafdRY
c9v099U0OZvo68oHxm/iV7hTp0qddz+sewGYG/Jp31mTdWi09Nb2MhTYz6bf4hvIKjq1DEq7CuG6
ZlNeKEZOguUFI7gjUaTpRldkRiLk2phiHIzS+A3Ans4d2CIH+11/GlagJ9xPefmDXU0WgWblnjFt
NAeErUwCj/aj7h5rhKqb+p2i09AXZHl0TxgU6M1xvzwi4Jr/Tva26snOOpL4YmRPp1Ix2OS6ATdm
ygFjBRSSuB/hSgFjqfjJG3e4P7NE3NUWQ1E3jSi+OBwwTEbSUixLrpkd+UTs9qpBd4hdXSPMKLI6
ZZwGp09L+6baw/NzHSg/7tZGxhfDtoq1Rlu85UpyJ9Dt6VeA+MHdImLIIqn+jxCAl85vST8ZdyZT
1IwalxhNkCr6YadpXuVzxXclcOlHU3iBNDXhc78DU3o92+pk6uhPoJ3YN/pxqCCCrClVe1J5WWtx
x0Uyxze7P0SmpaAn/T21t3bT19hkSBwDe8nduKeBbBTvpu80zX2h+bLKIv6vWmBu81jOqmbH8rZP
ELMzV0HqQxV2g2J4qCgE/EAf/lDcRgCutXuYL00Jz0yE93NCnMSk5SDwE0fKqL7cfruvAOgbSvEL
eJlSpWaR8lB2n6PnwX1bXlBSp0IJM8Yqk9eHEQl3UTDkSUlmzm8yrz6GNWQ2K8KMLj+UQ+mEAlXm
LGmV0ZjrQdTCRfoEKLSZZ/3GK4ZJLYp2Wk9Zm0SgLR6sB4ont0PgkgCxve6N4AgKpfURHwIitFyZ
7BhI0D36Ju//YTgLy8EVdsGKgZVWrNGK8tl7+yQlh8JGMP6i7TUH/HNbVdUwYqHZ8PEt61fqx6O+
90akyNgbXxxm7OkTx/HH2/oLpPa3kYqwjxfh25b2jQKNC8ea1G19TfRYHc7eOSyS3emGTXc9+GuM
6rqnmmKMfa9XnSQjjB0FT3Z3WBCbJp4eXJoLIErU5ohGAfF+FSiSCfizfvF+oENRfkkeX6KXtvP7
b1STmA+kKxcp7uBGGNWTEDSFtzuSajYd1jMNMBFf0dfLXY2Fl1bA5oacplDB7PLu9XBVWuwm84Kx
SkdiYknE4bJlTb0VkhP98UIu9XNr2nRpoElISUExu+AcL+s+Gx2vZMPYfyQ5N28G2wp/CCtI49lE
amwFSaiQOY7EsU76/CDgunsMn9F3ktYPwN8TOFFZM3Cb5RKeml9XRewC+1puer9WPo3HzYUQXWwr
+WQohTh3Z3dY2U0RWvXRzKfAFiHB8A2d42J0i9hCxB/tlYWxXsRuVl0E7B/1ZkEDD2jzhsFsZwZ3
IlALOE4wOEB4aYnC3NDYhcr4VEk1AZX/EI+6s+GRe4XdssIeJRPFBl/MK/6noQBZe7kIotozz+7P
eOCCdSczCAK6rhChgK/kHiXhYBiEvIpyWfnK4RkqJtkMxGGNOfIwFUeycxfpWUBfXDaImfOJ/Ua9
Q+tOuMzs5gfyk1ihqI8nBTXEOFBHZqLLtO4WgHmw5LX4DL/PkrH7i8qx917PJs/1uzle91nAsInB
Wgv89KD2XSSSiZ53jz2gLCKIPn6Y0ihDIVmkRgg9hJwsYz2jNmpcCUepV6U4vK32c8edmR2b9M3u
UZaGHfG3Vdfj8uAm7GesaMw5oGLl0uLBd3JXt3pLPxr493+pdqLrjGdS/JXZW3x1F0vTl/HVBZYy
8PUdCQk4lZGlUSdu8IS0StwPk+mlxnwzva9sTYMZfk3ASRBQIdWLcpnIJek87STl0an0eVtYg6Sf
hV2z9Z8nZjdiiq7e664E/JW8uotgnV+EQlmIcc4BYd/qrGfih5PZDKdoBQxnhJC/HKvsldD6cdV6
yJ8QEVr37UfZgUgWOnMh6G0RdzIo/2chWVlJkWDcy7kBjLJmvv/mY7Ttx0a89ncmjxPy74lcfJzG
TPZwegB74ixHdik0cvr/845iVXgVYuGQ+osgAx5hZenwxwSgLONEsZCx7MpjJe6TSCsFP4ygPeQI
hLevtfTxfBHRqJvBbIANfNmCWEC/SETOH1onaKw0yAxjxQmxHkkOuGg9tTSueYmGYg56Hr9rdrGn
gPi7nGMe5cbxZThsDueMTg8F74yz+1gADqVw1SCgmj1kuoCBUPQ2OXuCiCDj4fL9OWo311unQjcl
3TQ/VtrEcEH7hRsd7eavOTQw5oOcJ5AoaMQMSbIszcfAlcsQXgfOYa3J4c0uqsZ7/7tJRKorT45P
9N/Tq1SYD89gT1/YKNoNlpRlESepcSdmbHUQGTkOnxE0JNLnsuAJwPk50lFR8PJTl1GowzHVle51
TBzABW1Lro9aX2r0Hrf8iV4kD8GeettHLKI33HnqrMWkatmqDvHlYlZ2bd6wfD87+xkiCaaWN0mw
0cKKQOFz2MLRv6I71pFzWjJg0TWxetb4UcTqr1/UtNAqRI9OhT+/DTsAJftwfZza+U1GKr3vmQhb
iLT4WYlQqo7qIFssjTKMfVzh9zDj1VwhTrd6liEPk6nACFIH8Di0oj66/DCEY5dFn9HqpCnD1Zf6
kxlT3HNeKwPbeZjNuvhmo2r+Qxy0Q23jVHm/+3ptH2L8O5hlndQYZ24IaAw2w5vV6o38L/8BhsqG
GdpndYr8RTuuKmZBx5oEzjS23A7Bog9ODj6rzedXIILLotNfmRk6ZPDErlHr4aHs75cw5c8ytIpD
NRWaiw2kgXVmBDtmwv3UaKZmH0iF51usD+GglEM0rsLZUgSPilobSqfZ0KwroLpzgNIG6NBuKXGH
lDEWeMFxcPMkkAEHNChoihkf7Ui9/MRASbNJ9TtuU1jcgFiqUOS/C/wnnsF2a7zenBTfLFJJWq+I
K6LpdqFTH6YcbWwCsERjYr8iZTHo9KxYhsSsuB0DUAuHdNyiY0hwwaFHbv6UI+ctIETbsTGu6tRE
UUOvmhudgrMja4TzQCsaNqt4iBdsjaX3eAsUDfuNhDoqiPjHFYSsQJVz9yw1oOeB3A8vbaVDXs2N
xIpK3y+zpQ8D3RXCSPNvKJKIeYsljaQnLzCxJ4KnfDLxZV5WIVSsS4MnZqsbUKfK4g7NXUn1BVh5
cebFuptvjlBGlq4aWeKGSesQOnhAzS8mRo8QI0PX+5bTgRxnR9xUDYtfrtxueHrU4pfl+mSanYPC
se74i5VDqBSfvV4rzv7dZvICY6GmDLCCxeGzKHGIrpdteE8QCRElJEwsoKtfTToO1CS4Xv6Q4S9w
Ze5vYbFiBdqkDGIvgDZJ84CWvkmA33zcP92umswEsMcdigqb46oUqNNpiFOb6W35e/8tAQWYz9LX
+9Dy+3FUDCpZv8dNEzbK2xCPSn5u37CTDTdLN6wUDH+lv1m4g/lzp5Q8qpdcFHEOI/uMtdvpAX1q
z+0puJ9mW0LGDTOnpJqHprDGFIWWqO1QuJaA0K97xE5vc38SNwh+2FcvwNEJn1fLs9WqT5wJfpY9
obGplHW3X9Cl3w6FSymwPKGv0Yb8S6qwv+d1r8At2XYAbbpGU3KWwf2aL4Oj22ZVxdY6/gVS51BL
N7JudEhYiUrpHbziBEo5wQhw/hEGtUymLY9keOTEAco0N+cFjMpiJur3w5DPMvhHfXbneoEpo/hB
z3YMtKjDqNWreCHzMZeCto2V7maUNu4spITHDOBhL18G11SN4J3Dnsyg1WJIs45mKASFxNWy1bfq
cEgOV5hD0LWSDm7SOSub6qcW55yGdQs5FQRW14tAZCalC6HGM4D+wb/5oCcsir6LxKpRDlGK7QhG
TXw+Lawo70MQyB9y7v7PTJGi0ByLihIOYrvYvsLqFznhzrQGJz2Fd8oydTN5EUQr5jk2Yn0qCO2u
2w4NIkh+9Zlw+VqFZLXVwwoM/bucA+PWzga+ya0PrGOubezw+VwJjgMyIzxKJZmkAJkRFZIvqhH8
sat5mGqsSmYcgIHoABkUXbp0jnzNahXSqle6a5PEpSXTB3uu34LRC/dp1vlDi8Aw0kDQIfcWk2JF
gPotN2B7xUjiKy1MmMdeomaeKi6pGW1poZhIL6xxtm9eu7nQT8TNP6+kY2gZmRhtQc31rUPn4KhR
LY1o2lLpXpp8TPOrxKxkyOdYNSSGX1FunZRxDh+s8HX6FNbv7OPN05unMtrxqXKP8R4Fcs464Sp0
VJyU750UMBqHbPpRz89koKhHb+zBKUbNtMtSVmMoXadTHwri0mZGL1PrzLuOPt/U2cwGAglXlALs
mtuO8E+B0qPMpfHA+7V4H80NGMqoAhq1hhfOgNWvxyASsDZGvmK3X+/OR0LOUvparhrrjZGK2tVu
tVtsWoLDoSiDkeQE9a8GP/bJFagauwK9n1llECeHZEsY86agqlHFAQUza56oD5ospxo9IhuXUVJ6
KcVILXDi7pjdofZVs/1UcWL3l/Hkpm1EniE2ZR1K7M5Tzf9536gta6dN92vEq82WVRmdAMVBOpgA
NAOijKY/FEC5I/BWHrcwdSMbWGiBYahQfvQcvlZiM6cjFlKo/7ocV89BDEWxxBe7kFmoRhmfjrnN
OcX5NFbgdtB+5LOtND7iOhCdcVbhV0tGrYv4LKopXFkJmWFD7a65yBxqAEoTL7bHnCyyrNSwDPJo
+nk3DJGJBg12MLn23ldaUfcnbTYlKxEvYmuKn8nrhQAZ2hy6HZFpXSc/tE3Axbp74SDQ9z3g0v2Z
V4Rui6qQfwjZKlAmrkR9og9kvWBGbUNC3pSALDD7DmMi7dtE733wjGZ/WIGxWI0eifTeMYBBa0zQ
tNbOPmTenF3UmxwowXAMDU4GBOrGB4e2ZHFIw/d+W7EHK1IwTd5VW9f2y8p1mms9o1uzo+efv+J0
8TU/M+SGN5fy3q4Oph9aIsvOexNoJPe1GlgGl0WbDM4pMxsKt1nbaeQqvn1JAk/l/tsIaMstuBT5
YhAWd3yMZ4iUWKqz2ftMDTPIIT0rtCu2g7mexqQ3Q0S9uhJmwoSIudZBLdW4wGI0ycZnZ5S/n046
be7C1TAM9PbuV2lfiOSTSLngfmG6ajsvfKtJ/mYsgEya0mFgXf6uqXF+PXhic/8GLn0C+lQl3fM8
xSZMzgO7qHYFfwB/QqUpghS2A9xTUXbQsyx30Zw5tbd69g5IDhwygydbutki2iugbZmEw8w2b5FP
p9+2ytQQYbSXSqBhoxn2tLYjCJge1ywG4YtQYhVwC+hPzgt3QpciRm9KJXm0y6+aaf2pl9pUS8xo
4BCPkc8HrU4dhCAfgSzA4mzoVv3GEsdATIoUCRTnxF0XuCeY1d1iGF99yg+mwLlFr4eOzD/7Zl8G
MOsNKAjXmvHzx0Aoo6FsaOJz7gZqfHp+S4L06NMEJD83whicbt8YAPjTFX+km5jv3uSxtr9VxguY
xLAqmRUUlbLcW1pb7bcSIU0oIuxPlAyw3xFYViNwuvsiiIDCybuo06aVeISmAIlcECVEVApdGVzZ
NdKXWi4nGavmRxrgXJIduvAe58syaeYGUeSQnHdKwbXml2Fkd1bTLgktfwmzccQm2QNYoDfikqD7
F3htrHHEsqf6QggFqINUswLBONGtmUWVZwPwmqzKbeGUSH0Hn4bG55pI4VmXIugdZQnLXNsXgsHY
GGVBqXQjLaAP8eNEBvI0S6mqZholWOIll1ozxXNluFQRa7M78QBeiHDcZ58jOEtbgqMfLCWuAqp4
sXjECeTchWQepMNUJy4Q9nEQ310MD+rmBKjMaYYZ1cd6kgz5RuByXOR4OyL0CanEOOkUUgzHHBd6
fgsPp6QPAC+RUUZoxHXY/e2Z2ZJu3IbTWTyj2COtw7Gh9m/gqSirBTTzAv/2fsYL3rcQrV9VQFEA
w2tQ6n1oE770QMjjhWPyL0gOvWD7AhsGMV3Mqi3fR5neEFlOaxSnchqU4/1gR6AzkRx/pluNLboS
+hzPd57OfHKZ1MlfeCfZX3/Ck/vlykd41AKhmk32ukJ0bwYhuZ7HjvHTeZvIyTPu2wyklxynx9QW
DoT1eiCwjJQdKw3wTPe1tBCFRDywtXjqNsMnaUY1WG3YFHh1vhiaa+mNn/k+8sMeydAMfB6SUm8W
QPjG0wKrfBwv4uAKNR+3OtijJnnw/vDhyZ45se1Dk8XYcjlDx+zpMgokHQ0OyLr53TMoXl0aIwQg
9gFRG5AwNfUfVcy1ifKK3JEaTTeJeDWREhE9pVkETkw/DxXMIsEdeQ/sXrNRT5RYRvj6GNt9IUjJ
UBvNRIL4DAhxz2mbeUvFT8Hclu3YnnRG4/k3G8M55NoRXHoQ8RUEIpAynGwM1TvcB/dTXwp5o4KZ
60CpBWIJqEFh92fCQHo5PeN1bWE+LuSiXf6LtmHV0Xs6x/N0rAZ8gXWToD3+z6ujMzo7GP0kfka8
Oyl4GbrcknZmKj81FMBvATXmbpDRog1b1sI6+sZHrrV0F0n8275xjfVLV2ZdG4UOhOjLk5eZ3wa5
W5UV8KNN6vXUUy0Vm3yNCrviIJhlW1ctl49PCnNuQI97yATPtj+G+OSvINCFDdIHCDyRdqE2aiGa
JaJi0E6c92TWxTySTcAvcKFqMGn6U8WuHabuaes7JuAPj7S9bOuCDHDMp6mXp5epG9clwh3XyOSr
vrVp6OwVqC5il96X3WTjbcCTKAVY/jHKzqPHoJdzygz4Vdl2yXXbI+wP/KFLphLgy4lErgtocegh
RHZaf9DnJyXHrZzjdcaTO7GghGLcEk49ZemhRSCmTzVc9EYAO1kB7CLVxbOW+87h9Q4TNENKFr+g
ei5aEFZnEX4j8hjIW+BOzxv3KAGLc0iv79vNlLrEfp7VHPle/uqrYngSO8/YGTCk1W5sdV+m49J2
VPtruvYI7e1yDc1s5OghQ9bpIsyr/WSoIBFYMlXhnR2WMkPLhcWgVynfL85ElmJ9f8Vc8GoGvw5X
yq+E/xS9lyel1lo2cJk0t42uZ2KHkPstNTuWRIYro7+GQAQKX9jvuonuLuXb+mDMm86LBcwngBQl
aggxCPv749ILeX7hhAC4vSzOh/nYXNTQPd1mbP7IRkXPA6LpLnJL1SyJ1pCqXzW/dMa720QPwZX7
0NiFHyCW7p2/1xe6U9ks0HJlOZ9KGhoeBGCtBIKEWQLdnmIZEj9VNYT98RDofBxnWBxBo4kRJ/3j
3nHrbZrMY04hkKVAwyXbA0nkAo0x1IG+DNVa9p8Z26vLAX0mLO7Osa4j2CIbpAjD/+yy0ZM23sCz
Q6hWTeEpo5AOhkebXD8WCwtPcvegbIMDb8s3Om1r/4gJoLrqYkwWGJxJZVBG3xhgISMA52gp52v7
n6YXQ5EeqeEJdND+M5JyLQJDVoc6TeYQDX3ZgcajIisVRNcm77/4btABwoFJLS+QHS0h8D//RCGz
QMQMrhlaRqZfoQm6qkytHTjmJ1vESd8/XkaAE9abV2KLzgimknHjh1uVTwbxD4UsgCNK+ceYyapc
rUhEx8vaztt+BuURExNMyiDiZxIiF4VeJ2zTxLNh2L1E/KTew5MkNEyqYWLGG+W/plWg+IrgF8DK
eL9GHpTbekLcJXMBAX+k1CSaAZI/9MFRXib6Tmd3WkcrvoisDELKdgsu1YENGQL6oyJNDyMRVG6E
DZZcu3RPAAFtGF0zesGIwxmGC0B4chP118nOHBT7OsJRQVXRCvZsDSKHBCzXuUToEbQrG14vo1eX
je4P3A+Fz4fc/yzwGfuJoDxuuIbqjxmbCxrdCBsr0Ftr9lsT6aDGLVj5y8H8KKRshuI3txo/5rmQ
93kVszvOTAGZfFm2XpJIO5yGRWcmFhetRMPi5Zwx9y/89hdrvKeo2bekQobPvxta/Qlx8ibwQ31m
pBObgJhR2i+pMCD9OcP7biKkD4RPbxOFIAaBtuAT+1dz/iRImiJINqOMq3kfYUx42s9EQjgiow6G
V3M9ZNChikJ/supFU/i0ODCrfRPtipONM2fuKLf9MInUb79eisABLmUkzxUWB3/rI8IIBnVJROLu
2DBob22o6BdkMGYkkxEnQtIfVWbG0Jmgizw9VOBveNKE7ni8vggBjTXjOIk+LEFQ/MPCN+JKzh3H
p+xdiEvtSCzL1RuFup8Z7UX5cluGqFX1ZUElUl5LAPRTBdsTZI9I7Av89/4cupaws/lvuO6mxPSd
nEXmecVz+wj9TLOeEMLyzBcUYkYlFru5ei438rCEM1Y0/jwAJPFGptxQTFuTRgIIWZaYg16fsdGn
RaZ4mml8uATT9cshRuFp42tWGASxDVxu5cs5hp9GcwHwe3zOJNwiUonZYYXN1X9RhvmmG3mcfR4a
0ezrJ1q6xWddasX27ptyeT2yb0/BcaKK54bUlwube1Yd88GNjdjYRnyeALfsWqQMAOJ7ZVHDLIif
sdn1HWOSu5WvisIKeTJrRH3mHILpaDRB6yw1l53FrVaDeMUjZ7bT8eKQOfg7pm/zKPK7Oe4rntAg
YZkzeZ//VP0OxDRYFba9DGeDd/i+ACSjVpvm46fTnc+Ll+0Is6rvTsLzDVI9uijOYbEmh8gLBn3i
NTFSwK9exL9Ol5dDTR+uN6OTScx5I7YOkhI/OF7OZoaUAnvfDLJlLTJz4r/prS85Uul3M7vYgPri
okhnfcxUdYeIOwBCMY9tN0MtwmNFRjkIjRrTcvgQO9lbc4rpZFnBR5azMiHCBlFAAqm95D5WVeX9
Spfj0FYLBYHTW3k/ZPSkwRpQkb8PKF+ALtXMUHshU13kcgwzMk5Nqvq2I41fy+tbkFEGbtMm9LoE
M/hgmEI/yTX+5JCsMvnI8R7qTlhTmHVD5XbIubn+Uhi65Mvc+mvvtuUFdGKq49OmtDYNmQ7npHlq
kotO8BXg9g9tafzTiahSBdLheTHZpZLlh39AQdpcgHWyA32RyDWGfIXDwbv+I3aJPMIs7laKPUM0
/EpZ+3BwEk7N4xSRfl97MBfLTJTCTMNt+eZAW+Y4aDelmnfmkuQBeXNAIs/pmVWK6MuMFLxY5uXR
Hwzovp05ACvr538RqTn2qKb0fcyx08MJUj3/HQtrlpN5AHGGOK2uWFjS4DErnrOlYECd5bO51R38
IbTfklquVDZrEm5xo6agifZV4x2aRZUUfXWsbiZJ4+cVDAysAvu37a1xsHYToSwhXQPRLtQ0OsfC
7rIoF2z0fvNMoSZxjHB4lhc8ZYPlGW9L28YAuK/eV6ZluESr0/Qm381figu8nKfBn6cpmo2/EgXf
vA3XjmF3Vq9G98pWVsBq2eRAub2EblCqnfdA47E2bkSpiZ3Eptyl7LxlRzbeJVCPITtL+8k1+wOf
pgHV46uQ+fHwuoojeibb4CwsPjWOidY6PXUuSEGBcdxs+srRYcJIYdSdz7TmA9svglrLDz7axJ6w
U8AlorKmXNBqZMcbLHExYn500r2Jzi0/CrFv8To9qUrgtyygDx3/GeyOQA6FrymOv2KXLnSV4n0H
nW9Xv0WAhkP0cDioWYXfbm2zOEvCGtinT0P97hC4dwGDIZyYDb3WC1Hpnd87oc/zCVfdRtR58YHl
v5wvzfPkJHhPIaVdP8gRAjZ0UGWSeTJGKtt2dy71nK4ystqy1rL1qspM++F2U4KPTF+Cj9VOAQlq
80nEkelJnvMuUH5Xs/jE/yOxzLl5HAFDyXi36+75sRI4CCezyqIuPtyWRqe+iIM68R8LyIVTiCI1
hRtxwVa4LzuKX2cRVrs3NtfJWvD3tGBMWZeQjS52G+7Zzvu6QEHnyPNQ5HCipUvqAXu/NWZfOBxO
uKclF7CRjwuvoEFQ4OlUhFNSBbub3pTPmctTsndNOe6y7KnBfwixeKfAhrgsJE2KeDwuWWifHOGw
7O0w/S2DGw7XGC38ddbKWxj7Wvg8iIg2wrWtMWHRAU2RA3RD98XXgCb2D1HUz6DrtszzkHiFyMZX
LFIVuU2SXVeB7icwaQdTNsAzqL2+f8IkmzcQnDk5pxoBLwJEeb9Dv8oJyQrI4NxJtCxrZZvBJ2bW
WAVqGA+Wfqhcm096V2RBEDqGIKNUg/UlPhUQ3Oo8I7Cf2vwxRel4RIPlaN2cgSQgKKoy01ZKdY/b
4DDaSKWc1g1OGuYunf7pPw7+r31BH8+dQDTvhG7Q6BYW1UdbtBQnc/w1ww0TV1tFxOyCCI6Rxhyv
urXkX7EglHV/N5UdYQ/46oC5PagcRxvWDQ+NEsbeHxnUu0r03EjtYK/cP/K+UQogKwATaOV3wEtn
E4gYzrIq4QXQQ53KRAEJPsVAEYaJNULycruWuUMUjJUbj8LtEIHS83TstgPGdzbqUjbOBEj/0kOq
ZIUrnyer/SX8JqwqYKZY4m2u1JXIGCCwZeJ62/BQy3dmtbizYCnXAxPndSKP0l7/z+GVF8sfr9h9
bsZIE8u1uwy2QqgMngxVztbwhoYN4vv3kyMhq0zKjE3HpTshhV9VWN/yBk/4ar6ScKYGgeFF2b1x
vXAOW/zrCIgzshmTYBUBpRMkN27RuSxOXBzC4wgcS9QiIuHBqvXdQYrfj93Ei0lm1N3nAsJc9zDM
1kzXhK3jKs0wwdelBoHWMmCsK2mNVpbFxAFWMEZov3Pyy3Xh0iUQdln7BaAtOVQsAcna9gHL1l23
+XAdmmpeBrgSs9gWYe/8qdQAlEyuNr6yu5SOdH3nCAGHykrE9D/Hkt/JfUuPGjXTAczAqYbPRnGS
RUu0gIxo8xZkNJyrFG+BjceJxr04ia0WrslCnPZ/724UQoOsC9dCO8oWfBmVNleOYix80fMWR2xY
XofBBSoLfFK4nEz67dcbwmuIhlHj360/x2l5xP/SCx8jPB8+/8V0KBSxfuxsLOihz3x4Oifhfb0C
cKDPoA2aDDGvM5/KzoFWcgDBy0GqOLxoaCdy8CQA8AQF4qVqmcJ9DbVc/NS1XuLOrl7JABWJUsk5
i+k3EWnHLqoVirIarycEjN3aYb5lIKTCvI7Dc3ovji4q5IBLHDWSIvHk63fLbAgdf0w1sZfRQRpi
yczHKWSJQxe3Bhz99JSYewoARDwmja80l/vCQiXaD08rupGbUn6VOAtboE2+q14sSp6aU/1N4+wY
+yVxO6ZYuvG8DDrSKSBQC8DImYfY4EoXQqNxC30f5oU3S1+JA3n1KafJ5uameGJA1O9FCLZh9/AK
womXX89V7vJCggwDGAdRBy92PQ/x/xvupPQBimgU19lAGTBgHG7ixfs5nMEGQj+1wdEtiUh4Nt1i
e+c+GeGumcONN8yxYsLWAufMKa2TnruvcO35k5RnxVqFEftB60Zk6cttIwORAleWmkE4cThFX5kz
XpxVZsurSy2EpUA1NvEv86Bkar+AQJS3ugt4RwXXYsSxnAsyo+RbQuXuuX+C9fXtNurXSQo3Lw+D
3AezmeE6fHCnfGA/m+05y85jnv4OEG63Atcja34myqw8w8zfpFHyWPgLHLkfdtXF6Xved2YvmXUW
t6LNCTcv1OaPuvuTHT1HYUKpW3Hc32B7wvm+8Ww+sfYv3Cy1WSAL56Ds0j9NPDouR7pQaZQ4DeH/
vGZgWCblpXlrvQ4eL7KRUc+ST/5cDHv7HlAJnOyAmqGdCBMP58ISW5Q8dVNujCW2HikQrp3AOLIS
mlu409A33ow7/7XFNYrOQ3uy3r8piTnZDlwIBtfMxhE6h20avuP3IofC9BbJHO3iKI0CrA5sB2ew
sZWhU4A8XwI8Sjk1p6Awaou7tCBju+7vf0oENRtYrNnOQDX5aRENkej8JkSkQoEoD+XMyOQaGH5M
+7JDllZ18nRY2eTQfxqC9noYZLWSryay5Jq+Ul5G7lnGYw4I5sNnSypCVyTJ8B+j4bt4Je+ocHhi
D7j4UTR8bUZ2yqA4felYw8clZqqGgJmMmko=
`protect end_protected
