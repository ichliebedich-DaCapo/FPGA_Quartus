-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
npcK9hGNGJF5/aVB40afX5iP13N8DnKl+2fRfOi+78dtrDSDWCQz1hKcYFuRm0blUYjfeN7nPykq
6/8yJQpjUAJrwMDReVGrk8pKQ8dA5Smf/0bfUVEm/uCzNBIfxatpIBlCciFPS4N2Dfl0DJUedGN0
YgsjYQZ6qi24zYfeMj5wHE4c7KtW5ymKwnEJR/WNcaShpJF6OTaQMTVyL1MMep44IEor0Iz6CMQm
RlhGjMJ2lvyw1HFqeNHmOIYyQJYx35jToYYWBJvReUeWAMmycyoThpZ+M3ty9SbGkydneMXHHjLO
RPiWce7/VDum2KCaimUVw2HPWsrLulnO9LAQqw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14240)
`protect data_block
pKP8TS1tmDzAlH5CUQqmVAzRr7ovfTMk8w6fp2cMwhEQIEbzdFBEuiYjdv7hsU1bJ4YAuhV6PFna
U8Yyy6uRRDY2MOJNAwhlohXRpoIlj9uWlbcPc35CD7hK7T0NQz2u3pgSokjtNkawQpnlvT1EoTjn
qN3baOIA3oRoINfJK18rK1n7FHyODtF3CQ6zioyn6Tac9skjlhj192p7RIILvXxEg0spn/l1jy2/
4Od8LUhJ45InQOG+r877pJBSeib79ePrZbm5eePnJOdaVtk1acWEt5HeqcG+U+8qSOcSWsm1ECzy
0mHKHnTPVBLAUVUedCbMKNOJTH5v50R4YqVSapWw6oyUWCkUUCi+uENR0o8qM+PzmCKmpRqh/dTy
6QfGVXFaLEvcSr1JfQNqfdrMWt5UpN43+//xW+GEZi7GQqlGmhQjn9/R8LLcfF3M3yy/Fgf8PSaC
GL2y5FgbzboLopbyM7BYn02SpmOqljNud6pCinyADqOOo3CKCfgaFMmFhEhMU0CGDon3h2CFHSpi
ikPPvckcvgoKDF3ExqV0KHvcDC2CznYcQNhvrh9KVAtiDguGttwoS0aJqO3jMPWR1LdqFC8z+Mlx
Ry73ia0CNLI71z8BU5eDPU08C/7IHZZi+MsXCxuaJTFEuA2QF2AnVLw6iyBsL0mVw0bOzZgEx08R
k81CufDtQW+ADh6sJZh4DZPqYsWmTOJVJ832k6j8cVbcKWm06scrbq5os/bPdEXUlTt4InB36VFq
rGamo5EWEPvPeISspi2S4pxL8x+qka/UNpq369OSjwCaGtfloUQjVVQQY88p+GZ1FFyHDNDw2ip4
nUz9rkmzm+sffBL84wOsasY+yb9md0yovX4A7JgWvf6YCnAJRLpeyvkHMK8OPIEdNe5Oef6rR6lK
fkejasozDIBvjZvzO3wxHNS8ra+bDRuibFACVm2L6pWWPPaAV2xh5oKH9xfIA+X9yBeQ3t+8lMQp
Z0ksjKbPjshPA6Y75sWL0JLRxHtm0l/BzqEyEDE6K5utB18eubviw+wvnZGFal3oyS0hUQskLRju
i157vZJharO6ZVUJcb2zdHn4o9EpEeZyPKlvILCPOg3UG4TCByC1eVpWEPMZIkerGS+q0DRtJaid
pvm5yMq4yQ/iyG/GUDk3P04a+fv0sfvyM5oUI9gtZsyvhjrmIVoA2LxBjC+VqQQHxOWk40mrac6D
vZbEKVZaqHacrwl1vDf2cBSxQJRmXvGYYhY7sJMpd60dgEzcdn0JMCKjIIMH5t8zX+AK+41IaU9D
kv2mTxQ0br8oc2aIfFu5IC1T/c+ZNe5W/b5+Ocj95KyJSLQ4QglAbKU5ySLopqB7rEJk+43s8flg
455c0Ne6rd/1zgQg0lSG91HS8svBlMYihItstfFyagYb/va/PFsZkuzhE+PXmOR5CcoVk+ml5Iow
r1Ugmi7GyKjJ9LuQPvZlfz1AFwm7NI127Tdu9j6D4Wb3IHDXbVdFbM/XMLXiXzk7+5x9pFOuLIKS
OE8+6Xn6W2iUl09ejjgAupgiaCIe1Px2Y0MkrvNVk9pAFM+Mg5hVfjwt9Z8K9i1MEnPRiaVm2ZuG
ZBt/nhNk2PL2/68+hDoCbZgufBHn0KOTFaRJ9zffn3uSfIZMX0+IRt94otTDwRQfjo2jcMJZXILB
rdKUlVKl63/yTi/RzW83OaIxESb8p6xf4PL2Q1trZ+uq4I2N49Emnw35jUwwjIn9lCTZlcr7aihW
0Kg893hes9KP8Ve+c0Q6Xgx3ZOQiRfnpl0pMPJExK4rll/9PSxrQvqzJ2R4j1uPzL7lOd2hRoMAU
S+RaSweDExivkweUul7I7/f5CboxjbNbjNNFXFeVFrFyiHt4RAtQH7vpjHLihLHpwYRlqyslz6Xd
pCNOa52hlrTGhcw1lqRl2pJ45KIwAeBC0+jbEciu3v+hZAfyJCBOOyf2QQ6xPlPYRDS7RiWSix5P
Kf4ULMHvUT/YJua9CY6ZJe/YQjL3yc/IAYRQvdHxfSPIv/DZe1X7y/uuTRhJ9PqdHT9bLoTa7T3G
ek7qqAYP/W7lH9ue5AaknIZ3T1raX3E6beF3SclkhNrAE94fHOx/1x072w/X997m48jj8El+35xC
sv1pomeLA7hj+gO9tu/fg8MBDwHdiKa5rmNu5iAiUHIb5YMvFU1vvziO/zfMP/tdcKu2tsZghO+p
+ZKhOuZ/zFK+l9I9NBpfpG22VzZs+4TU5StjodldqAd+j7L3JO9w1W3eLBj+wdADr+dPQxl3Hygt
VJl628viVit7hxlVGnkCqcqLiwuw3TCNKup4Fdk1fWo3qdYWwQJ7jdR+woP173DA8umDNMbERG4V
aCBP9s27ieWZfH/uhccTKkHsSpYd68ZuNmYqOLC2GqD/eKeKvqbM+tIfmDUX+3djq0zBKalzBNW1
Ch2FUfUHn5J8Uth8F+jSa41uYbQe+deA/dZJcBZv/ncckt72XmWDe2OP4opEiM1HgTUQOVGlFrGs
a7Do/BM9AsX1W61/L8ITk/cFo2wcyhPr+sLZo+ERcOW/bodV55yIXHSgXR6jBKvpmCw3GSxy1R0d
k5aX/nQpyBKNvo9Jr5K90jL1SqJYgBsT74KjkLtV8ij9xyFWJPK9Riogc/gPtvBtBNj7VCflLj17
a2Ak4k9QYcQJn7nEZMLGGgE6hEwgpCnLbkko/aMvrtTS8U2BoWwW7+c+1wNZjO4RaVq5mQdSdJBh
/Tkf3jMyS6VljA0mIA6Cv7p7edqK1zp8B4+cCwpnCqRpu/Py6WOt4pAMdXVN9De+G1Ga8BlRaqEe
Nyd1X6NbfCFFgcxdrKy8tbMTAOXswF2IwMaL/9XLlrcPstdcy1DZNw0TKq4kzOkHZIV1UAv5kX+z
CrV6PlVHUVGy8D2inn6pCFwqmIzOKt4Kb86zS1oCTusd7Px5rAVaPAQ3KsF/cMIbBYCEntfm1P8X
D/5lLW4Rbi2RxxiLMpoLKhi5GP33xHCctXLAW9JCggVSzFqbS9H0ce1w3Jw2xJ+ZTzCxXGpW6yVy
vPdlRAY5ZHsesbTKKpKl4I8SutwzEme6PHqRB22BNnkkqaeKh1Y2s06HKB2m8MSYwSpFG0VXWfP8
SXjwQi+VD8c/LawUU/W+6m3fsE1KLm9lCgQZ0peQgMfInn1xOlLBrdxIgi222SSqsJo7splOAJm+
8ossL8YFCwIlaAXkYgTf+2mbWb6p2VFn9kyI3TxLG0OgCYcvdAStPPwaWetjAtZJTwqHiKEHl16O
x6SQpjtY5NtDWSYHqTTI7ghxMdm71/7f+ngew8M2b4oLD7QtE/o9GuNc5+KfO5vsMLgFU3AApWcz
dOrJQK+2p54DQAPZxAmussxLvZlicJ9Cpe6v8aNGdNsz7ogDLVo+I3xNRHwFT5L0/WrOWenJ/MkM
hzsUjcr2+9cksYX+EYGTkke7sSYUVI1At7w2IIuteGqkbRWiuTyf71dEE9wbkOIFdOC8Qc2XbY93
j48qk6umQUDEhPIWC31G2afCiG17lIQIizmjuJ0XIwhXzzQFFANG1KPGnz1wDErRwpoWMjP4fQru
XCOOrhYegj+5qotw1fw4Zs8O7Vpvmy1jf7ggJ2npsDsO9nnVdwOcZ6vhzZVo7/hF7UP/ruCCgzcq
Ioz6hY06juWYYRxqCVimijgrbq/RZuGFi7H/pTw31s7qogbOjMuyqkkgNlcaMejR6gF6S8NTknOt
2i8e1EJhgsR08B2es6zGyMS4vUrb1q4ni4F9hSWX2PjKvBZJ8D2VVQMTbcE0qnhAx7QT4oGyEY+H
+6U8P6/ZbCE3DKt/yfJeeQXlfRSC459cZKNGQqgkQJhzYzNduQf9VTVwTg0upA+JYNq8PD/YgPNt
oxrBa/gF6jmjCudkCHWPRzmXEfoPDGDPFiNLNgpRDSOZ5vQ4BIh9uMIiW8drrRfMli3l07TbLg5t
Irfnr35EoY4Fm/tUrNxWB1ip/L5J6TITIrNs9QFB+Al7huflyfOE4cgA3sZZe3GMd5lVdHWOygMy
Km76qC+JLbM5gqjuAZ3V9S06G8lMALu7tTUW3HefLZRP/8CuyHpqmt3Gxr4/X0NyCcP2q/VhXBAw
5Ty5k2OuMv3I0CPYxj7NjQLPktxKMEb7WL93L4PMpTZOQzGZp/b90/hg/xczD2K4ZJKvr8YLb9rg
wXrz6vdUg59S1EI5CIqLTKU3GMJfTpoKRoPpOFCYQB9Z62m10TsN2XHZQrk/0cZvnm1LuFFwzmmE
sjWL0e8v4HcKas1Mp5soN0GVpKufgREMWrx8zKUCEbEuxpjd0pMJfQU2NpbezKIyASBjRoQWBTKH
tV09/01a6Pd2XPiaVV1czSLhGr4zreTcfc/Pik4QtqPI2x8ZpeFLtITdJBuL7LPPSK1eANQG2Imc
R7RRb7BaV4doN6np0Nqhx1V4jYtWCk/0EN8HqwzoB8iAUZmN/bN3b1Dy2iYQTeuvBTa9mrRIQDID
uZ/0K/hhlyFba55th5APS2AO/4dyBpm2/M8G1HNFkSlbgzvw5ByfsNTGM7emeeMqeySHwbQmJ6wl
PvkwMGzRUjgDMn0E3S+7twR8/DoPKf1zhb2I02j7UhWUtPT5Vg3DEGcnTXRE++CDO9PDXOwQq94k
NC08aJyKbxpgrgkEg47IYeH57J4sTMbhyYEaKGp4KaiotHMBxi6UJifPiOsWqAMuGL3ewtGtrAG1
A20LfYaLMXnrVFTgpg0JVD10LVpXSelHMgmcpv5l2Y8JkIJpXzobFDgrNJzVSb1O0MKjEdigUBq7
dd0aS8AuxpqHeXfoV5bKWtqIJ6Sa21FUI3nq/TAB10HGtbuD15Vff0fPzdfhh80dZkuX/YSmCKcF
WOZy/D1zkNi3jGWnuhzlOOdrd0oQg1YPf0y6SpFr6KNEfOHJUcdzNy7AodXE/ut0svgpGs4yrGLI
Eg6OjC2Sl6cGlbwBm+N3HL9ynNP+C89A76yPbmpsMc+M9oML8kaSgkAtoUHhXh8PSdwYr+Z2zrKc
pNIc7uwelo3qwbq3HLi5byZX6N7cLRVlb4NDC8D266gj6f1Xxd/yqJmzgIJU5enbamZ7L81nnbkK
TNcOBTxV1Q5IF2kwE3NNjE5e6slN2uQddzF7yYQoLlRf6RweIeqIpfpFxk3ABcMHB4848+oDL03y
t5bV9doaaP5eVkqLNzGFqLe0A6FA50sw41fX9Ug/gmA3PXKm2LQvcTPtJcXiq9u8XD84yU9FzGzL
wg6IIKp9El0tTgsqCVeKI9zWw7RH0P4dgIxpG4zL8D8yE1TXbHa/jrRNcecB/lm8M8oCfeDxpCf+
KXX9NPsXOzyAXB0VlCJAbVFCZDZadFQiW2dLYAH8EukilDK17VgfXZuqL1wvLsxzXbCQpigZxe3H
FtTvwWyS/KodfyTI5qMFdNKYfzoEOxBVDVPDmKzom7NMmQNUMKK8IcAGeASAeE+D8Q0pDw2NTkDn
gCal39rkTO5LRkxGnRvDtH5CCVixNcfLQ8a6X+6uJNnxQ9XzhVzQVgc7GXLpmjhJr2yRb7mVol0k
cprcFqP+HR1QmlBvB0KXmVpCVNXszqgX9AEljTtbaUICvdJNr7OK8N+Si8K58IciUonDlTQKdPlK
mpzBay/71jAMAGuBFWBlv0vhbB8kENYhtESo9NrlgGAERJbuWa0+MXascEFkaqJatQ1fA4/mNSEL
m2m0UDsy2TJ40Uh1bGUgwUm6d8WskSnKgA4rrjQs87bs70IcdooGADRXOfUd9Jl3vLvfWZezUWfS
lyH7gJZ+6MK10D3K1I92XxNgjj667uT/WIHczbQbHmosWvqTAxuDo4eVwLt+OUHqBdHz+K+O5b7h
aC/cgKwQ+i8FbzDbkTAaqc6mj2Ltd7EgPtrrpo3dCpgMKntIYnHNku+spouzKc7U1J+61Uu0MTpZ
DKQ6q452ET7dz06donvMvRi0EJSFYp13aMmWrqCcoGyEGqP2b1vNfNTk2e75BJG2KuWhHm/0lkk1
LXY/zsCdxm0Wpu4tmw2XJ9BsUn4fTWEGjScqtWrxweNZobhiOWFZEYIxS3E9Laj6BMj+f+JLTwIL
d3Hgurx9r5D9RMcbNsYXxF2dkO+W2HYGd3Ajg1L3cnKNQuvzjfB1e4Uoh3ooCyFpp2hQTRVCuQwQ
iE9AIWxJ9e721I2zgkwvCpXfujJfJAAgt1z1M74Fzo9hSU8d2UFy4O7YHr+CPRPCdo/NARLY06uj
BDS4Z5ugsTLdT7ME+1/LdXixVtV0ZPTcldmqHvoxdiGabzTC8NHEsqCm7kt5HWrKx61lWVxUlQam
QNFUeFHMiXCOH/qrkRSWArL2V0CidgsptHxdzx04N7lfT6tfdsoBsAR5NowDtRBxKo94/j7vMSpW
fkcCzXkQlOXZFvUK3/MLuUAprx2M1//EeiYYCdfmiVe+MV3vg3uUWEmBdnwYB+4ev3A2ZgIm8nuK
Yur+cLlb9S87aCosrgqUotnrqbrlre6dPbu0s7F0UsCQTlIvTkGXlBUGIU9pOxShhX0G+vv9ERm9
lcCzWaZWdM4AZ++ZB98qEEY49Ln89/a0ln148QNvkuA9358PtOp8dQ830L0ZOHim4U9RXkpnWog+
1jjTxo9O/kiDKcMwQRMgnyP8L52pCS5+0v2NQH2Zi33YBGif/CGfB/CIq0jF1BtnoPXyxsX0fJHe
61UNQ3JLeyyLTTC3tvF6ISDnqFWmcw01bWWf6TOhwkzV0lrmN8wmIFVcIM1AnR36vxHkeOgNy9uZ
sPA6OwbdOjth+PfLUaCmbE6k0l9Rgepb1sKlC+W6ousKlDyKm50WqNwjgSHjoCGRh/mu7X8S1Rqk
CtDraHQ98JdcI7Dw910iG/4hqfXkhYnpA6SNsYqYNRiSZ/yl6vodS2YykO40l42q3ay2ThTg92mD
55vX0thET2fVF4pLEHRIugNKr/oQTdIva7JoPmEzodKg726HfVMuz3XYk4RLZ/N95mcC9slHyZx6
erImZBVLRi7i/3OMYsA8egu4+9CY+n6u2P4/0HUNLXJa86C2oQe5wQbW6p6Vtg1BgqxxlpqEHozh
/w9QCvlZyf4MW0xqvxJfCy17qgK2JrFpMjiA6XWrnVc0AJG8O7Jk9F+lo5QxCY/tzHYKDkbO0DY1
IEXTzrQOs2PkyF7XnhWUCjJiPcLnJevasZ5AfgTYJucvwRkyq4+IIEbDBfcRsiCwacQ8QEMC+RFU
0haPEuPs3B+QvfhLGgtQCXgyTxd9A+xy1a+mWJZG2L8nnuMmq+up+rmveRUTxpPDXqLQRxCZCjOx
HWskvQJ7JUKaPzT2302+lK0eAfJC14aG2QX9e0+VQ9XKJrTUKB/4laadmRoHozbDhKN0i1jsYLap
Lx3xO0hhN322bI9+gRFE2L/Bkok6aP3NToQylWUwFMZ7PgwGWSdqjFB9kUPhLJ8bFsE4/FOdXzRl
SHOoFJhDzr0lkN5I2BnPjEOuI212as71WESvpV5AebLpEjK8GwoWXmJNHMPr9ygECyIBOT4c6r9c
fKUAPquRiYBUsOfZ9CfcO/8uHSJxjLTyguj3k7TFBhERWoxGVjPrvTHh64KI8JozE3ZrVFmsZBkb
6NIFNXik34LngSF+XnGScCsg/7fVUVTOn96Qo4HdbY32WrkXGLbtNd8Z/pti1KmATEQg8rVprBKS
XpMT1+ilGDltJWhRFO0Qhhuon2OlfF+Z95UHZF/ef8aMf7+Ae+Lrp6FB7gTMpSSthieclKlQOdKH
W8vkdkT3HeiXHdWw7pMnUc318fLPyqZ2RldrTxf7mxtwXB2I+rKRSXzHXLkui7xrJdwVbifAxbDj
f6t5fdza3WzKU7Rs7MGyGUWSxaqVRptBeZtJ1h1aD8XRpQcG9iYtU7vUXJkXFpH8xqRr1EXiyUok
Y44fVY6J4emMTGtkUmn7z+BYzwmd61tNtvBVCtSHj1hkpL3billhMVFZejLoQqVR5vojc/Vdie1A
Wtb1Pxmnei1b9DwJUZd7GjJzYjoImg6n5IYFcVSlyx/PH0S5sZcMtR1zfLsOMZY4E6wu4hvYvJgV
EmhaTT0Uw7x0Vo275vsA8bi0ZM0oEHm/9GEaz04e93gokyKinznI0c3HF0QvdtKW3wWWbu0u9Hfq
+d0ZV+1dGXaRCgiLMzVQC/6VpPMAtqCq0Eey8iPMMJJoG7WwxZzCBsg+CTVsF+3kuKcalkDYo0Kg
aD5KTlUE8i4V7XTlRx+xbzPpbRvVJoKwHDhzK1oj04cL+Kbha8A7Gx314BZb4+WqEmgZTUdaUxgc
9fqbSPQYBlxFZoWDoi8rPI4woLH+VGk0CPmmJoZbhMmcEOfKklFueGAvwfVmIQhLhgUNhrBpEgtk
TwNzrvM3nytH/gKk9A+c/7VycTsAp6xpQ81LBXrd+eSXuKwezM4VrahU691v8Fw7guNq8Um9HYRw
unrAgamIeoFxLU58nBO0suhsN0Ba4ElIUy4wgaTlYPrP2dyOyeQbtWhij5QZHOIuKnTUjF6rNCdR
YVKknDPByl9n499fBQH204upcjkGx2C5hoiN8HBYKDlDQNWNU7yf8/d+k8Yz+Yvmowuj/CWdqXZG
JtPbPCsNOF4K3vxP81r1C18xS/auZ7udhtmpWLPfjrfIF+guN7x1oep/zdDkfn03Cxp9yh/EnuCe
f+8BAjh83x0kymvr6oDF1bL+1pnSvwxNIOa73LwU21CXegCF36Rk2Gpg6iLUCxWigr6tEtg7RBYj
LZw8iZAqVqfM7q0Q96Fym+iZ+Bn6cAsFOnRjv+3UgAAcVEjrShFCM8dkHcyOqWkISL4q0ArqrPRg
EsY3e5DDQi7f36hexaY0dByXNibUoC48hrrhU3y+QBJzTWderjEaiY2B0gpCaOtvYHDQ8vKhUpme
UU3ESoFOypktyG1jqHL662n2/jcwvJ5MePP3Olrv+9CQ5s/M7y5Psqv6AFe4YPsd+mhniu+08QrU
y2olBBjLivbvX5mDglwD9SPG9JFUdDLB+CirA+TOsKOPbPXEz/Re39einekE9mO7HSw+YHTmg+K/
yMGKYybLpszf2pK1JQr/vy9U6PFkqu6gtRL/wIMKwE6mO37nxq4gswLsrKKAkYsSN27rXz7VtRiZ
NgspSy9JRlYy688f0n7RcUvyMbEOmB5uX1Qz9n4AF1/5y7X0IYhjZwsIHOOSfBtc4Vw4Hg3Gk+aO
4tMsh06IzScEWMzflSmEe/ptTKadwuDp7DTNwDi6AUwJT/s6jne7Xd19z161cM7aC7hVbfi/3dZ5
3rvc08XrKtDGTttZg3uNl04/msJVdyBQdvzCCLHH3H8QxPZKaMfWi/OJrVQxrC8MDgI4So0w5KcH
TRGlUx4HBHxRUklRKONmXUXF+6uMsl7iQe7XeK80VGPhzqR67vEuw1kQAGDC6dEsQ6a+gxUDT5lV
VeaqoHJbf+B/WmW2at7kXPKEb1IwCKOCxxHXaa7QSpC+kBHn39G/Ak4WTB35XKho4Mhpsst2YdFi
ygKTIcApX1Hzqaps6oMuHa/IoDS6QpZM7NIEcM8lefYuZbGhsGUyVvjxz2NEsh6nM185dk9l7q7D
N8bPnuWx6wxLm+FlCJW/u2Vq5mOpgViqn8GvAV8uQ2V2jJNuZImQvavi0arga5Plx2KATEVRLBLe
fa4fI1yGBFyPkHBQ79KSE1ssy2JsMFz65fr4OeAL441AfXD675HUByasbFpApYlPD6G99NWSmUKL
u+FLdGdhvSkqRRw3NmcKtLgB4/bJ1WVEkshIFt3nE69UwVXBWK7ZOi94NCB2GSbNqMcTB3NokcBq
u1LJLawTXJGXVvPd+8eme/lDyxBd/9si0JLxdnMxijI0pSXysyaExItwhACoAm6BjHCSkZOliR5O
i+Q2Xixga2iWSUTdKFMSRAiwhATujCXAoh1PWgaQr3CsJMBE4tN+8iaeUHWpOSgkye79CnMXy17B
hgjk7RWTYWT9cGrDOpVqcL24g+Grwc3MEGDE+I3FXg2sZk+kXP5Dooj8Ktkjeaf5REmltHR6U4Ud
/30Vw/pCMaq2mLpoipJVrA0WbvXsJGcl4cuKq7WKM5Tvw4fP/Y44u1+uNpSSpSRsYn1IQbfAJXYU
ROB9tM1NESWj8ZuGR5qHknsJHq150qxwiNzsSE4IbKghty2tsNFrLdruvBdhnlU8EvcEs3xNu2mh
NNPXVkk4/0FKqQ5k4UQc5BbF1nhtVm0BdXwTk1YnIOkjbp7hiRBZ7woyHLAa4COEC9HWiOwYiW1L
eU2g25vQfC5xcUAZpwlMGjiBYtqMxn52aRdYW5Z2BwDYFMYHNPpuQiQ6z+6x2xUg3bjKt2geHAgt
+svWywe/3XYY+VAXktv6ILWMXRmdF7p0Ox4Mlh+PzK3VEj6gY3sIZt01zpn6IFXlAmdD6tsfvc5N
J/VcfyWK4PDiTgyAs6wReETmozFGLbvY9AwABQM2dEQ81g2Z1yquTM4TTwKzJmiPWQCISsBJU503
AFjF1k4oScPTj7131gcqYhMVRDgRlhmcXhTFGXegp5PGIfU1GbhuZjCuXE1HrPvzd5peY6HvJ12F
y0+QXUdYCTP6PPud8+fRy+v4c+v5Wnd50al+NstA4BvDgP3QoJjaNF0EC5vCsZdUCZUVcyoHurMi
i8e2RyVk6fNuE5Wt2ls3ddqMvGnQBNQOrvPLBCldqZi0o1IJKdIg4cpRHpCGPxMmgqsaq7z8FIwC
/I3HbE++spx9XR2ebB73Oq4VQHEjNABmsU1FiRmmw2aL6VcxKb5hYtrgcFoPhqzIyYgJgAPnAVnQ
zTOryzOb0xXdDQfVPYvfciS0rSh1aZv2gJ7ZHxqs7tQUMdK+ip3Iehsr+xPcM1vgzmjz7LpYpxs4
MLJ67tCruzcobyVdlRqMXKPM/cqhHneab2Hlsw364ieUw/ZLeVeO5yvODh9zDw6lTZEf+EJp0kxx
KxStxB3qd/TSXFV2l5CkNIzr8wKkPbDheyhbV4pCPLHBRNAzgAKCmoA71N688SdKu5HCsEXPFdYd
4W1jii8A8HJHeDymfxHuUPZ3M1eiAyYrJOtNIjM2zHkXeuk7uQ1Ch2JA+JXMLutAQchQtWy4fy+2
iPd8Zmp/bjehqixEtuS5u1ji8ujzuJIgZJMKRspuf6eZzLD6Ua5fHD7Wyel48xF+XdtHok3Vnvj5
3KRMg+ZFIVIBWeufSAX9yA9xCHov5ANmA9s9OTtYIBUAkx5IL5MPCZPc0kc9M/L4ZowCiZ/Q8qQf
2S02sAgjnDTrCUzAKJJGbB7+KWChihLlMTGb6XhP/kOVpaIS4s4U/y0LuvEg1H0XLHY342Ln8sF5
GXG+fwxCeIj9f3zSA6KkRZSZoKP94ZaQI6DqLXvgxEw8ul89k4Z64gtNmFZFYHJKgBiPgl/CwUJi
9lu8KZk6aynNyTn2QFfJp/DmSP3WS+GFP9ajF3TF/zdPGMqm9OaihtTEREFUxB5k+6H7aayXBbt/
woir2ErqjVpWpZzjD6ZmRjASl0PnoVOa9ujL0lYKBsJXo+XSBzjL+fjbbyCz/Qyk1jBfBP9YMjmL
mWriBwWHRkXm8wrOikdZWCenr6bfm8J3pRDeJnPwkiDTHrKAa9u2jlPrMlhEHFz0y/znMSHm2qFj
LiPesJoZxHNvklypl1hTuQFlYe/X1h9eZ5OA9AlXiSISheQk0Pxu0GBvx52g2remyRkqJfV3iS1N
2Zd4CbpjH6ROvJFqyO4T8aAMJucQ0xYU8DlSxcABU1t3D8RPyh7hogHDjKUPQ9g0148JjMZRzJos
sV7oxWGqI2bGGNm/BcizfbulLgaDORtmJ8y/YJEYzAX5eg+NXBuZcPTrpgKeviiT9fw5VswKbV1i
iNWJrC8CquubTYCMtQE3Z5zEQYZmazU1803m+4+N0mxPNSVgXrbCQezHc5o5kvMQejIPeaiQ1BQt
H5G318zX01msl1PaB2vkS/98/bUxrHv4BTsNbGSIk5Jf14ol2cqRhCbsmz3fXIPQ6D2yS5BTvXH9
9Jgv/qG7++JzzDTpl4/b0HqZ/vj7oC0SPRBe7xUDbCi9S8F1WJ08ZbxgsS/it7jElvVSIBWN4CKG
+EE1fOxWwNbY2aHRlSin/dhc6mWFu4YlS4pj8szHYQuY6N3Tn6JEwH7oMokW8HuwMBKHJQ2MuKXe
LAYkFXNXRe9zB0LRuWCWo0Zclke73p0VbzQDSYoS9D76AlD4Ahbdc6HhVBTc7OpUn1g1emXpVUye
9bzcRhvlL645hkNPfRvTvPCdTc3/uCX5JjwEA+xMNJxtgR5EaJtGzJZQKsn9l2MkA2cbpiQ9Z5aS
3S+IlDQ3HmWnNeZyE+RLHY96cemuLz2rJ80/h1aUvRSysXQqhQJJ9A69lF7nbjgbSM3ONoQ5S48G
FTJfFPNpoN2juTB5UZnn39SMxlkksDov2mw6HPpSCoVGGgz/YqwDXUNTfBqCF4OfHpELgGg3rORW
07QEvNWo7nvgfnKcz5gsz4QbvTx01GDwW02Ad6Mvtj96G7KUsbz054svvBwJwiEwCsRMNSlCHkbS
NRzLNVnY1eZW4Ir2G5gkfh7k5TSaybO1xHwpM9hKHnfbmUkKyIDgOIH98UwgUby56s0BbRg9EWXy
FICex8+PVaBpzJTZuTIehy4oJBFo1om9qufJCQbih7F1xI1ENNr7nIcEuqpe8uD0eK1ALeGwJ/sj
/Qvco/GxbEpa6usZ+saeVI/kNFK1SRbTKMvhyA0TTmdYk+HP3b4b/tcvQE4qnFmXPMacWYph0hho
1ZRxyHx1yghFaIL9XKlMojySTVTVUNAQ6hM7Ly9Dk7ka6Bdbhfv2l9LEWQ06ZgDCXD4EidQEdmx7
ac5CGj0sZC/La8ej9EPsNbVcpEhd42/S/DH0tMgnGJ7AKvsDYsjSa6M4ha8F088v7eaYBcQXHDdR
5ehEkoF8X7O5YckXSOBkpbE8E1aZRyj9ZcDhD8CoUA1HHc4ccr3BCy/+mo4Sds7ViEbv0Lh7XQZU
/Eqxk50g1TKzSWNC/zYboKtqaO+su/O/pz1OPJZ4vGSf9imTSTlg4qfYrElBb7g8oaRae4YEr6EM
Yv2PFZut3gCEmYDav879OkRkTKjrjCSVvfZOcIt/NntQnSYeCw5kYy9wgHjMByo0k52KRIysn6Dz
4TmyqLnEKFkvxfeTpMHHKFwauUrQwzgNpUAMYV8A3suCOe2vWuRFQoWFxwR2Ciw1G3+bgmmAKr9e
qiF3PEnL4Cxfjt2Yt0d+BDvqNrpvPjzjLTMo5Q9dyHlimUfO2byQfUOkS9HAIP4cTDBteFc9xMvS
m6KBRZcK3a68cBNiLWIQo/Whg3K4I/jbyAO+fACJFrbElRw/nn7mq9DBnyecbeIBa830ADDTCdnt
+6mkqdTKFzceupf8xRpQyTO4td64tmPCQRTZRekoOj12TFJ3mBPq/besvicwvtrO6OszJVptT4GT
4d6A2GF9UXsMrVwCvJDXHRscSLwAcEokhqT0afg7GwiuItIv9yjUDH30FbgY8updp/10R1EesBPf
Lw7fLpK4luDEKyyXdGEBo25RM0Yp4E7swf75DM+C3AYD8DcxJzoRUOmqYR+eDRrWddpc2HwiJO0x
nB13JU9oPcXccYrH9zfdc3/NHUR6uYYGOKGDqtXRKKYOMZw+3vdx/DQUkNrnObq2ViyO8Z2Z5/9G
LrIW4kGg1S/xtUVaOj9wL7Gz8WqdunzICS6W9wJkPx4p3H6F7D7wMlP9Tz+oGu+NRXV6sVuV1Tvo
VkT75UGV9DG5r/FErQy398tzHaMVZD9UdiJSBeSQTK8jQZeDWu+MTH1AmHN5Ec591HNhHIrMzBif
eD+sb1tKTs7CHQzXgyOnrTpZhxQBY3HT/7IPEcd9ukoEkZBHRHXR/g4UX4CNh1JSuCQBeloRmcG5
qNL2zu+5wnrzFY9NMcGtfHs/TTWJc9HDFpcSqh13OfVp+I8V0rjyEMEmQZlg81jHV+13wWIwNadD
UQ4z6dY9VAr6GNUi1ClZVjp+OggJ+yVmH9ceQXKVHDGFkYUu90D5pqLeeDbHP7OlqbJdaJhUPVJD
7CPU3VgylItjSVYdffA4kl6Yy43JQx/9LLSU4juak3qrgjbK7Sbs3FdjijhG9TdEFqWrqUTO3tKP
+y0aZQrwM1iwH1Fw6vmEP4WqXikqZuv8VhGaGeoZt8/tarCT80ilJIasAwrBbQahc5OgEY6NSFs/
C29Yb/W92P4Wo3WfUqPMXKR1jwJSAy/fZdSaI+7X+ywjYkdmV3UP1jXlG727usQyqUESnz262qZa
efkYDviuR/eQHUaci92dkjLJ33Jw7UnMtTp0xBZ/EAzHAb84rraIMvMRpYkNfZGdBKntkCRvSgeY
8YNdVo4Pb/C/OyVefIAMrGAhpjo5N80BmEHhP108hBM4r0eB6SAC5m2u6R5yHBYy7ijn1NW0KjaJ
y2xDsCSWeViw4nH10yHSVmK09z5XOKQhNFACEAPrnMzvswsgiY2KVsDFcTUhYbpGOg1bBSrBuvz4
YtpcgjjYhe2YtYM2dhKt9dU2QATCiQXmrxbi2xBOnVjRNUugCd9n+tLNDIHKpElyBe4fv7rX4ryt
5+fdoQplt4A37TcbSiOkVK3Q8QCvhjs2d+U6wBPtV7c52TYWMOc41wLlM62vO+r2/4GN1KH279Nv
4V2SrPcZ2LkGEymjk9tDq/DhyEvQEwdq3loLpB3cMB5e0xwrSFoGPFuBD8In0cwh1YJzY65KTEhi
tFCwHAkJt6OVdT1HdGmcrTvsptCY8cc3HA7rU4n+eu57XS18mt/t+ihmlLKMTbZmXj19xlKiXyvI
dIC7zCVfDT29s9hb5ERW2Uq7fU5Gu1RTZ+9VVo+CeF1C351MyVoDXX39ad/yrmSKaa7Jr37KlTw2
KiXUk1yn9GK+De+5GEVPHg3+nN32VDkT2ILkiZcPAM3hBl+eqpVvca1Si+qWoV08jxseB/KI5SED
blTzu1cZE+Q/K8Epee8NUHqb3CHzm7ZLdd2+aOYSnwYuVtjDOuTUgsWimYGt5602UH387Y28xMmG
4TM0n1KTnBWE9J/teqppZSfKut12/Gi306qR1clh2tdIkeHqO5KMteeX9tcnKC1zrEDSSfy7r0k4
qTOOJr/sI1IURxWr/5kXwbzn54EYCb3rE5/sO/1j7XIbWo3KU0OBKUVCqG6JMhACkRtJH1YEVot1
jZCmP52hkea8DggoryxPzPX9O0kgnQEqjbWM2KZKwvaUlE6aCtej5q0HTmA+STTjzzm95wDx4eeQ
AlETgR0KoZUMZPnv5zv3jm2e+PvDIffsfd+M9QqbyOlfiMWhwzntmLs5oFhbk7EKQvFURoa1I3Ph
E9sr/CLf5uwmLfUN39lcbocQBIR7joZElTgTAwPPPrtSVykRR7WL5HaNMIw1oVJTjsR2AieaL7/R
sYH8fMFfpP64gd7VfSx2hQqOgMaOv1XG+SUN/5a6ZwWxN2ylDp1Nwo8Z2UYH1vuRYaQc27Ls/1+R
KsWvxQE+xhMXwPlpFNLm9xoHXslvAIFZ6LD03OUfgzVbaLxCX/6tf+Z+a4oQFwtBL8wYnhLgpemx
ZYcccRTelEnry/rr8lR1HJL8ZesLPJtqpVATbskeLAu0zg60qv+0Uh1sUDQoY+VmZbq+Lz1WsWYS
m6Tc89R1jFJ8uWP+XbZeiqQG0IBn3oyieA4qJbRM6epIeStYigHnbdOX93Emd6Ce4bXukK0ts6iq
oRxn2mS6fkb/Qle9aS0sFA0574g9hqHMU3CnZ+ipS4T/62tAczZa/Gm25g6llv9tfPdPOf1AOYU2
r34INcYei9/gMP/ItDdoDm8oxt5d64TnfhS1Uk9JNaK8Ma0Fqee1vDMPKreoMhjTSXWkHUxiWNwX
lswFOaroegW88xm8FwQUYO9dlxYC9wohGVuG8yr33Xs3fHqn73Omq+6YLUmNkFbMGw4v/zhN8jho
0nEEf9DRjctTFwfUfSfqFb0FzoEeOatwHEYRi5KFxApJDE2k/kFMomYOHRg51armFKW/J2+/bpWJ
n5CedAf813Kl1UOVclYWKb44/PR4AOeChwCoMRdXRvBFOhBif12ZIuoCs8cUPnT88irxxEJ6zd7i
VdkQh9NxMpAJ7syAChAefXCHg11EbqqM+x6NSxLQYT0cXsgB7fFLZngNlgj5w761J65/DGlfpqLk
liB7rzfAzzha//C240UzOgG5CHm8hNBRalUjPZVCXy1J4VJx3XDWu1143gjCXwdi55cZyDBMKJMt
JgJguPijMtTCV9jW/ls9E4vf1g00lXhfqd07cclVtdw1cEuCcYKCh5L/PnVXppHgMJ4Bb75mqGe8
ChrwDHj8SDgxxMiN7V5sZOoLCqiVt7lPwNVeZ8BkoEDTuSv5nezTXeTGxWlHBAHeVm2bjz/uMVWa
K2YnxF7FbfgfKtwjQwjadvAWygpUUSjUuPgsm3Qt458CNXw+/SC/O0Wcwd1OP4i4/OCbTVtlyCyt
k172f3EQB/6o+Mp5KJ+43igrLGfy7aPeaDp+edeIBf4bzbDgoFvSeHcoy9fTjyW2sAup3yS1bh6b
REI4RkUWSwyyTq3E+A926AlQjcA/A0EjctsYdqgvWWSYHCKYWM5Wsk8n+dowVEGm6J4hdwCcQ3tG
pjFU7vzstTh2cnrwHD98TGWgxMAqnwEN8P9o1jga+Hq+PhY7QRlYm5OBAg5MobCnX7kgzYiIayjx
eV7QQlajTmosFJiovI/kdshQAPVJRQ3bGvzcJJbVXrrUoNhJKOR/pfNGTQqZ1PDocTneT7UMFUw0
rPGPEK3xV2mouJNC0pY6stULvKfk4gY2EiR59GJN6lUmLEQjxWdcQxmqL0WUlM7Qw8V2dgnihWlB
120jFGwW9VrkRUmcraFibAPiVUixc5J5W2Kc8Kxk1SOzzQAD7oLysvAJmshXrb81JsyK0T5rngMO
Bkw6bbpwfquaEkmqS3C9e3dvxqWtxQCbQHTpn97iagbDKt/tiXEHUqXwKkNFaIw5XwQfADVHQTA8
5z571dIUoN354BcrSpTwlzBzTWSItdmRSCVMyPIwlFqUucI5nUPgUQnWptLlOJR6ifn/LeT6KGyG
MmPPzTFcUq8tGRUargHqHYXh6XdXqHN0c4T19EQsRiC8O1Q3eDF5ZB8KAk0VRFlsSFNNuCJFnFZx
WR0DFA2Zi11lM/X2eVasOxjUwiYvz6fAN7ude5nFQfDckss+TpKLCN8OokHHCY4i5IGfUlcKXyfX
ZIOIEVOeUHKN/PX6FxtQ26rAigV1EUXhg6E0PMJiffb1yB2zY7eG8XfppvQsDoEDjv1HzAP1V/JU
amsrsk7qK/1I3Ms4tpnufy15eFNEsRgaKyMz/upei7Q8utco/uv0LrAfuwzgevLoSA6J49EZ6ylc
ZJ6yCzNhTYbt2G+fy0vKT+HSYagVgJG+EOua7+MdfotdyP9h/Ppe7veZmI2tGOQKiyENcOy8XfAH
+T8ZxvKx1iKiexzO1ezlAvOsdIWe54QLGx1meuKb8+cbnNDfb6QGIIYpamUFiBH4fOtJu+Ku/Bbx
VmUJmKS6mFSD+wvKslfEn5AWmfiN4Ga2GNTS0KOxRSDNATDVEnRBjOVB4JXXB+tcs5zWXTB4YBFI
TkNtZw4cq4CPEogVcFzpQvpu8iRVbYQz4laTrlhtimjpbFSDX5dxW/Uv0EY9zspiLWoSgMyGr6GY
NyAh+PUfyIOIfgc+wZERdKjWZNn5uxeBcod/K6YXISbnOyhLiJyoLjHHj1p35E7HQVMagn0puoQ+
DDvK3oiWdF9EhyeHdvKVdiepJgEioccyMR2pjgxkuHiBtQqH/Lv2ueG9TEtwYa4ejB/6/NPSfGdM
XK6ai8oGIJ0iBAVV/9+fVYU+pNvOcH1M/9af919o0WEF5oh/jaw5YG7FdBdjMHBMfk/ntnTf3vaT
VRDiBze0wzhBUxWBLEurczBXVKxhojvi6CEd0SxPUvU1a40B+7eVBIeo61E+oiB+DxgZ4580m8+t
xhGgoe9KqYIlZDO9STnZt88GK+AFNgG/FQeVR+ETWwjrzXNt9xhbOz3qLG7fUt/eGPHH3DXQhSeN
SHNNSKOGZLD3dDRCrkbAVaSeIzmOfKNTYPHqR9hbWiwn4kx1DZQkdAE7ktJ7xUqkjHUzrPtvBjaY
0/TNVSJ1E5C1nJ7xghiEiH5VdmemLqBSL25ioT6rF+sR/FvtxRfni1i7AtxZZ7VB/yMuAtmMtIeV
9IEn9C057rjgpWPjxe4Ux184xI3j/NbhUIS0gWEjhjNOIZCc8tRfd2Whd9XN+5UcEevm8Gdyyhtf
pMaC5/MpvW3O0N5VPGy06WvbypicutfpU8EHisJTAG543v38hl3x9Jy6P9WsqEXu/pUHoZsXih6h
8tjBdvdUpfZpaaOVbq0lQ3lnF8tRt5zVv3WCZBtmR+coVNjNyX01IT9H0lyzgKctjR7jh4nuto5q
oITT8ZWQvHCW5QlEMzVhq/kmUW/fiWsLBMOBWKIJJQ6Rvk3l0hs3gZGmBZwFHy8ks1Ijr6m3LvQB
LQ5pYFgSjZw0+oYQrQT6NaEi4MCbLUrmqdFaIYlJqK8eU4tUe4fbt01N/+/fwHZXctbAh1gyIbB4
ShIiMkudhpmoaDkYXabVoy7U0HcHhWm7yiHfZPRPZr+68GCLRiZLnzjg+5p51GKyS0P9sXD1i11x
Bq1Pgd1i7IXiqLUXnC4fhjT6YR3cVScf8CPKge3gl5s4LMKb4nX2UVWi0NLe51+tXIREsKrT7ZjW
sDxlzZvFABgsMVdfRWvS/XGvd70s/XfxYBYmtBkOojdXpqzvLotLJRa3DI3WnYNM5MNrhbhzLLxq
F+gK8rxe//Cny2EWsnTmqJ6o2gmG2RrSkDQKRzX6TcMR5tpN/UoqzRQ6YB8XHAEDn7teuEWmxJT8
mH46Yz4A+DTbS//+oNfngEWs8PdidvesgIVlMsMqTLF2uULOOvoYbFVkaseqkK8=
`protect end_protected
