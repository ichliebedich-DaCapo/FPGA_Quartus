-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DTTbXVeaOlMPWHJfXFZdSHu4fjhpWN5FApit6aPituyNImheONOfD40n9+zRQwMh6mpCz/495Q+r
FhuWUIf1Y1+FU2rklkLGDQT0lblJhIc2Bz35jvn85BtwXorG8aKXIGHqvTv4yhIdEkCgdxeGg93q
SVyIc9BhDY8pxuuSKTAYGJvrCfVHJjDGisvTR1o+DCw0DM1e1KGJuIbl8sAEWwBOn563sarAbZ41
1p2VArhRh+HRTAgrjCHdKvNToobT3P6fOWiFuA1ZZEQ+mkKy8xeY9qO1o7WamfE5is33a56d7hcR
QxRDID79QE9oLHFgosUHgVwM/j/4X/6QbmD/7g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6992)
`protect data_block
tRaXy/4cXe8Jz8WDqLdf3Li4FPVnpzXkqnTWDaXulWk+N2bw6DHkC1fnIpaB+GQLLe920ICWHa/+
JgX4WLqS3vhMZZnUsC+ZWHY4OM6EWbtRKhRyi2AUqw8MydkYAO/QoRwSPimoQ7OollSlVIOj7NVm
059JkD9vw9WT61fDiNt4RmEgg38YaQ5CVwKs4ahp5ocjTVoRDJROezJ4ckNaOe0OEyDin1gCDpd0
JpF0w/gqYg/zVDQYXXN/HJ02ObSLT3u83dr9bWo65LEJGUmIey41kSv9ijyWoDxl6M46Le+5Tf3L
sjnvs1Hep1OACa4RL7yE/xkJ0XusY6t+ThSILtSI8qqnKyHBbDTlIyrM6kvGLOgynSge1fMQs+Rr
+q+xmYM0zc31LHLjB5+S8C6I9GNvvbIEyiEZIJhmaurs/w0BXXBj6qludfB8FhmjRZKeAjORFIgp
vdVn6Am4TJB4FiiTkopvkGVShYE8ZPsS/vihW2wspVfV3ebZbzQ/Yh+jbeBLQT37sxF2sclqSoBR
m9VOIswDEoriW95GqvlKQCQNSk+YAoR9wV3k7qN3r+0zcqKLODsJxg7/WMMh5a7uW3h+n+n0sNIW
zI5xb0YGuoaI+vOPYrYoSuueBo0ewAblAqtwO561BMbaGK4JwqU3REwNjInt1hiBvTx/Q7/Qsn42
e57GvjIKtZQS/cqMLrtMFa83qOE2UfMxqmIQm6oaIubRd9lW92Fu+QOeOTqiPksQu1YqeETsTlV+
8Zqz7AO7cmrZGs98GsYS18VitBgRXRWXEmx6OCPuKc2RA9Ym9eE4LAMyrDqRkU7A1HNgXOLTAIRW
mlRF9DrFl3VmriHXNzaMO47oAi5+L7EkkmMI3bdXIaXJUFJCQsdFD7bzXazTy16LkOBto1jXOvRl
Wv0qGDqA9w6I+EQV+jCloy1Qs3danzrlv3CXgcwgOJmRIpEsuJ3p8uI7yBat6J0du6+1Hx1uLlcX
WwX82UKLmyeT01bZjghxXtkZQcj4QmTkqoPn3CslNvbjBc8rMWtX0A9osGZ8xVVB8kzofj6F8mp4
k+78IyFbRHys/fnvHOzmLC0fI3Ls8ag6FIeGYCST9gz+SXQqoYJOfgzwYDG6DaPkv6C+1EZt5/Kt
Oo0iXJFHXaS9TcQNY0z+9o7KMqQDX82AFxKjDFznKo2Fh5fIef5z7G6makhmgBmqZLIJezvg9pUu
U5vuUiRHbddFoHshN9v/Tq1PSalJrbkB89N8XidK+bngEBsp8HMUKl4gbz1r5o/HHHz94TNU1W9t
iPZ83VLT6roZTnpWFUufbkQbw8BKGKVuYTuOseme5/9AQ5wI+o9gYMKeabttFxbjY3VR6yb6QwZx
3P0sqg97qMQF/02Oo7NbK6qcApf8fzx/WFoPyBP1Q5ZqoZ6v3ofLVf2apTlmNMOeGyJzQLBhVOtY
rGpuA0gqWIUPKEmsNrE6ZxsCBcE/eDwwxYNgpCVCDKk0tROealbJCQfCDTlmRkBOuNvGlQLeDCJT
7103My58A8NVkkOuoetI3AUsqwXsY8qeUhgJm+GECHO7ejcR3dFcyCVFp/wleQkb6GRlY9Y4XrCY
Q3B90N0qtRFb29VgR+yl5JlYkCSY0pXOUyvxVMw+aOyiaYxyC6SMzThwvES9pT7rRO/4W0PmfKeK
NsNppLaBhm0QoaPSQzWPbhH8qAAKlucYf9TDj80eShMt6Yng1JU0rDOCHnK2+7vg0532h6jRw0mt
yYIg/w4dr7Ajifpp59l+prdMzNGC9GS0Egfe/nZGDEYcPIJk9ZFpcLMzReA9s6K66dhI0hpU8suP
1aik7jpHYpqH9yxq0B/DZzD7ep2JKk40APaPqVrJl23GpFacfAtH0EudcqObiL9fO+yd+CThW/Nt
bPR0eCwZeEC8iDwNeVRzWu/D099QJj70pBZNQKZeFvLFLafZpGzrnxUegnTHMFl8eSw+msmCfWv4
/RXFvk4PuJpKRfsBmxcXRev2nUVrtsFdkK1ZDkQOH3JptyTrzXY0m1xMlsIUwWnhiaE895qEo5j1
Cq9fM3F2k9Lfp1h3KK1M730WZO+YqFu1+fFURWQo5lvYY5gIr+vP/ayQmgjXLb6qo9CWZklCX/bn
GmIcz9iLazxTfa5tfpwMUDZy4tJ8AXBFMAKp6LlfQmU9oj9+BGUkXGoyizjTqwzQj/j0iDrmYoHT
Mg9cwAnlQWDJaa6uVBw1Ife/RRvMGvwZ10gHanrFNUv5bx25X/MpOlNkY01LYXiuB968E4uLWDGB
OT/GtLCdY/mexAYbIzbzfjq1wbMYLA9EKWrdWuftvvTsPmVNM3pF7HL7pCzZEEJALDUL7+2PhnQg
2QEAgCej7W3s8frVJQQ8Ixdk5GRNLkzmGwFTpeHvbnnQdLwZz2gxmKs9Ik9lT/FYX4NPWOL1l334
IeLTpLcNYdkmQA4ZOgqO5UmBHgwlZIrABXbzU6j14dL4BRX40OI1zCym+cCOmNqy25Oj6Qd2/P9J
Gl1db1SC74vmE0nLnx69NhqlS57fCT+cD3wVeRHpMDw+Rvk69WNpFYRmWop48v89LKpUccfxi2R5
jeGrtfJYEjMDkQJBz6otpN8pI7h7DMuY8HSlrQgHLULnysAgdTYy7htx2eh1/vLRz5m9zlygcl+w
ngNgvzToEqbWb0JSjTjp7pIc6ochHXveCXhiDPi6iU+IcORoNGFP+UEJi5bm/ZdVmKOuG17jssE6
niq+svk9SfM5qn3YFwRiqwSS+yIw7Kz2F2YjGBdbbNmC916FC7J4BwJc9YhHdW5fj620u9qMVkvP
St2+9AaN1STLX+iIiBgLkDyvayuqqOsd4rsJkYfc1xFToNgoKGpu8NU18garm4Scvp+xL+P4qeH0
0Gy06Qkz+Ci9XYO3k8ZVyUdKOARhYyiYI0idtX6NRRZ3KvSPVUU47mAXFPPhHgxxGWyMyVith8Sn
j+/G/GQQWgv0qny+iyLZYiZ9I87lyy9AenP4xIk9gItC+rVIhAH6rJxGxPOQN3gM6vchlEwg+KDE
87vjlS6+MPNHKTzzVHfNlsG6JDiPFpVCTQYyQMAURtMHvqUBkwKrs8Lepcx4GtnFiYOi8EVRsI8Y
8UxnYG4WtF7Sl8GED1e4BZ156fkNT9TIAv7qPe1J/QODAoj9ePSxbqbWj6vIv1cdrcREClYTgA2V
XyXz0UYUP6IwPooEx4cuA+MBZwYZJ6WpIqKJ0IyvznbF8SFxOaNZWjGe1xgMcZpJaOfFHU+ciQ/C
ektsNJ1DiEiKeO8QePN3wjkl9oEjh+vA7Ol9vaDvfohZzsBHLdEnGpmiT5wY1Ec+Syd2AN3/uGMW
hKQzhAE3Zwr2UW/5KNGGftPhXc3C10RNHd7lLLVAGDNPto1dJl3timP7OV4kFmdIQcptbp34cHgY
6QsEI7UM+il/ihaab2r6ET07g/L/4go83Bzq78AfzUTnzYiIk+TK5IcTwm73opa4vYNuwQQMXTC8
yE1pC+y5huSANyPpCrctBkYeb8fMtfXNy6EKxRepCE5UQ5xzgOsQWwLaHQWVJoa1FMYPj4QCkz+P
/WT7snfONMw7WFRnLU4BxbPb+bkM55TZ6XVEmnxgWZevMEFlEXFl/dV3K4B8UZf9ZgEaRZPey1Hu
/kCpjb+TKCG5ZESH4HUS0rIx/PTxKez7gG3AA0NyCd+UTTAGuKGMAw/2n8eBE3kk7jv3XNbq29gB
jAWHwyB9ralYWOWRkGSFvo8Rrwc89AHHgZqvQMCZWDPoW06asG3rFvzNOpbS+NsHSGkk0UoL2gAk
YeERa5mQc0jFjkO1jtMOzlfKLHZW5623IWSyscgPTXxaU2Bq+h48aJwGUVsks6hWTwdBbTRkBFhw
yM5QoahBTfslPUVAbccKp7iS0BfUxeMbTOXXgqbPszRv2uYMLODHJxfUc5RfcXyeVwSQLLtrWq+Z
lJhUJCrFDNuEn9OR4Ci7fVBuECj3alpJzqZ6lrySj/fgWxitYw9x9NRtSYNZHe4sMDPi2NTuiT+g
icUlbscJMeAonpWvyKCmj3kHGjy+HwAQDNmst+1qwvf/KdwsLK0k7MLmFYrjomogpWIBDstwip3d
G372wBjpDS41hOXSwQw2KAzqeK+CF/t0WP8lZZzR2B6POk4Z++J9Md7gQLo1ehQcnYYtmMlnIonG
0WYyJSs0wG7+C4ADtJlUHxaTuI3P1N0f4wCnRrFP7hXK59/l75modT4b3xz+9kifJzP5K2DcTYYD
nKrkPal0dkRP7OKCwrczeelQzWCe8hOZeHwByrjW2eHstTYusZJ1ONXuwSRUpLwUn5aNDwZvR04I
Bz/cKX6VQ2j78KSLFhXAnwrFEne+UBD6eWNUumFJpnChX4otGiZ4CqL91+q2oAy1XjhHE3wPtGFy
vIQujkeeVjeXjR/UbvFUWf93caSrkN0S/CyvVSYyeY4u109GqFp7xAHyjxAUbVSGSA87lWfpCDWc
99Gl6DEddmC2Ycq8xxCIaPRtAScHiHUSrce4raCiCivxKAX4E8v6NmZDyCriKD8hGjwOETjeMFRI
2dAzTx4DB2e81AqdqiNB1q+f7N9ilTJAZ6wxWFpY/cA91xyGYSxxfmt2XEYGYMQhqJxjR5KVYnWy
upqVr1N7Udu7JoJv9qqn3uO77Q1bW/3Bb/78W5M4mq5F6GygExOr1wStVEnNtCCQSB9pK99pWDwC
TD3Yc2enCU8jjOd2XvNhyUSrrbdPV6r1KbiKkmZuxkOfUQYvWzxJQzh7TSIP7V+21zPzjCZiWzwn
Je5QKK4Xn2lFOYZyR5/BFXJXh8HcgPduSiZwMVB3GGEavCILNaydtrHQ4ECFB07zGceTOYkSmRjK
hTp7OOTnIsR8+scu+z3SkAQ8g/4YL50AFHMvEo2oFdJmVFecXxNAmTtoV/V0WGQu6dsZIfWl2pcg
y9g8yDNFuVQZBMhrO0+jDhRC9aBowJMAztwmpqxHCXe113JXeXAELJJFBJL9PLLmHajHsj8fU+4r
3YEJNQIx+FWIy8OZMYn56BjxX3bFsuE8jcWVaCVAi0F5M+ShfKfJugoFJPe5JWHUuChlycpgCUPR
F9dc4llBAA0+11UxXq4uKlDNi2KtJ66BYhDObkgYC9kqG+b1EKz+6DzMVfc1o2M6E8OVz7syO0Sl
PcWDa1fLwOhSRTgeNX3itkcn0JN15iM5JR2Cp02n/c9N9QuJjFdanbeHKYKTbL2jnYnC/l1uLuEK
bZYDenHiVGpF0GZbluuu0HGHQNwz8CqoLZ4vyxD23dfq6Oo9KzL6LgvhDLWe0WCdthokONRq5uKp
wamZw8DzrA7KAYUPjJipkWgd+zW7za7ljrXjd9tcHOX3ih9RTK2KOhl/soGi643WLFFFC6vNEDqR
mUxbpeEW4xqSdOnBzGd5u+P3+vo7B06jtVPkdzuCRIMGdV1Sqb9/qhmdwC61QXVq11yDuhcxQQxf
1KIoOLvdsSP9pAwXkWYxFLOhX9gYyjr7zMs6MxiQJyyGRaqRkqmP+ngbtokIh1eHYEZfnEwBcyVa
5mdv/Jp5WrR/SwshWhl0wJMPjQ1e99Zo9a9VYz5pqNfR7UD7kz8F0s8CvCRCOuTS0o4amMH+OpXv
LIV6JfwB6iM4OTg43f1+GSI3vP13rp2DMW5/DJeK/Ht7fgwubaCoaAkFHZL4SDOW9qaD8KwyOwop
5BGPUKQd/MVtXh7cwmBLy/7HWKJt4GE1e/o0qHE2XkgBLg2lSZLwxF63CcqHbAksAsfUKHUfS/1n
hfOSC6lj3CY6RoIKrSw12Fu3hIS1u4AxkVaID1yDlLU+fWJjxHP4zgO7aiLgv9TWWIaCX7tiMTJc
72g07VWBxVvBmonL1i/IAM+J3m3Oa+j11VHJD/RnMocPLac5kKzXB92RiJ7oaAU9cr6HoXEnF22R
rinBxQTC9tyzxWVXGBV6NcvSdgnsgUkF6ruwnW9E2NAWFR6rXzeILVM37+Ele+slcfrcuFIJmJ0L
srR+Eb4RCuqwGPTmRQz/tFYLZ9kxCNdgqEwxGs3DvkzbGgJMtLOVpaKsDcSZE0UrtpwE4f5yWXFb
XDo9g2Z77d5RBRKcpXWPnWVbiROqiM2TmUhrBgY7KjNWUFMDNn3LqPdI/5icAwA2MgZ6vpPHOhDT
D6KNsZYYDfQAIMr1Tuk/nF3k3nWcH/PDQr+RHtP2/vw88yHBtRCvOtTo/wCkC5KkyJa9++dDdbdN
4k7IcVAldE0VTnip62fFtsScMqIEjQkalWyNM+AlvRZPjgkjri7ruPPmnSMtV/r803h2o6bfBgMW
kHw5P98XjVtJli6xKULwKV/hWjoL+5255hes9QXcMmU/DrsC8r0+dWcpRCgEpwkDoIfIUXMKdFGp
IjofMzBRAbJdrLr8JxuH4UHOfU9zTXRRVTnEPjJOIH+ZHZEJhRIrU20A9qCvKe2M8QEhgIFbteN9
jswrozfth/VordFGA8LIoA+FRCZlGRbf9C6eRgy/Is0iqjB2TJOvdqOwxCaxdAwDXU6YAjcPje5Z
eay09V3/tMfZ7rwnDVdSEBpzA0N2/dKoAvRXWB3ryZKLZmTZmiyrasV+Szb6T2iC4h+HLeKl7nIX
RwTo5VZBsLELXFQuVbI19byzTYWzVcIwRxNd+VvXb+M6NJVyO1NR4PxrrAXJAspEH5F69nBl4RG4
TFbvaIVfH6vw5NZVzgGNaWMFEQvhVkQJXapMa6pW2r7u8DDeaXQNTMAlLqsu2pbQYCVg0N+LZduC
Jb30LnsLOX4FUrzgmmeNdAKSIcGydZJ8/STVosvPT0zbbsXsZ5ZQWg6ZDRzsM/UUMNRZ/WaxuSlP
GVADt9pNc8jdxecq1d737jN1rsOyuJ6XED8n6JIZU9/9FcVPlSHSY8whQmIB0bXkScMP5sjPgRE6
Act8bPPM8lKBN8tp4/mqSu/soTYs5MxxTnZcNN9qNpXh/K9Kko/KqrR35bsf8LIdss71P7td3GAV
Ifs+urTWxHk+eht2h8M5aUmCnsD5Ysc0BudnBoJXlhVrSCOGQfWn6NWvv+qblYPYySZjFhYJ+OG0
XyJZprqYdBMJT9fsqwjmjjoOb7aFB6rq1ziLynAdJGzaYrRt/W+motAR2GJhX0HOEcnIqp8JY2Gq
EGpPOzioJFj8JoYE5ObyGp+mg3jvoW3oW2aflOm/zqm3TJHx7fiarLpcZFe6OCpj0B28NRnw2OhU
eThqzmnmpIU4wO0IkTeGpXukaKbZ2EhXCl6YP7OXzuLlEYpqSCEErRwNQmZnqvMdXEtU/8o6mbX+
bVH79FH2Dmjcu7VtZhPBO728CsgX8aD5JM5OcPNC8uqBmslLTqMq5WjdIzjL47GuS5bqi+cR25Y2
BtvhZIKJOMzV7z3rq1hd0QJb/Gqv+S4+45d+/YoSiqTJU5NxiahUeRi4VkJB0qazknR04s7A6Mgb
wB6Ac0jm9g57yTJP1cyr8vBlQC6TbEU6YhJ2Al/GcGYY2F3IKMu7aacbnWuACRF1h4WvkYKY/eis
iautJ4O1Tffl5KdeBEZhAUxKzCxWNzHbjcWa4TGZMzmiZhfm1h7pnFsS6x/57IxBz3b3Rnc6udZw
5xWqs+H0pyrZcVwsxMZRVXna9PdnbjEsmSFHQfvm+6b5lV+KtRql0vhmJq3RniL3LgLNs6TbgZJJ
a0ITYKQNGz8T47sXoKXB7ZhwzCOgQ98Qc14K5FfOjUggXMU9d4KsRgr9yF4DzfG5t/0I/VuAgvKD
41vOWdYxSvO8sd3WT8k7EOMk3r0t3o/nYy7Ynn8wJwQG1/34oF7xUa68FuyltUPNxo54kQ0xZcAX
bZ8YTZYXmdNk0K06bMWZSHem7ANLRXlTmUaJi4pyU+ldPQ1VSPWgLRnoouYh3SaN3c8WVPgwlNKO
8hh7CXuQiR06iR8ydhFUZ0jvQiSTFLZHpFRov7O8ddE5jGje3H4Y61hqrOlwQxOiEXCbi5i/XUGJ
MAhqCyb+AyFrhU3yEvnp+C6Tbk7uMcz3rTPEDYnClqlG4uQFVTjt9dmG7rm24QC2YCDWDMnqP/Yp
J3+FoYa/DIe4e+QUVOZ53opCw0Kvv8nAAGXMxP2VcLdUS70yQ30eGGrKJbUUICQU73vSvXuOIxf4
+VPUvsX2XZnLqcTxKoL/9VmJNULTLxKx4JvemVqds056yrysXCjzy8rVh2qiyS1OHsWzlmEk8xz5
aZSQUt/H1tmo//KmplWVNH8/BvEytbHsUcKq2dZEn7jNYD79usXKE9jRkQSXRsPIUOxBPS0Vr0xK
+Ksp0OWVJBgQgRha9YYAaH2eZ8uNco6YWw7oyJOImIVai3FhW/4a/XM1TFH/q+Nxq6kQufTGBvFp
ekrN5/nH/1yCmmuI3EsF5sK3zcU8nf87bCP0hpNyzzSrZR5T9GYJNOyX8ImBFfNqPy85EwCWEUPe
1VQ/zX78UM1/75zSUY9uOp6kH2NQBlf/WXhEjrvVOhQ3NHgAa+ocVk6g3dSuB9F5nyRBe5KEbNk3
QdaISZvdpcG2vcOvN8xRXwer38rUcrgKilRuVdRI7vGMzVMsg7+FYhGCBwTapjuw45TTYD95WaFI
s8fzJLzI/Vrkkyb0ZO9kKU9E8LTx/hQ8l3P/4x7MVzh8wabdl8ps1n76li75/NM1qQ9082BCmNUf
uIhj1i4FxkHO2cR8SV76NfD4tdkXRupvUWYgYmrp3pnvhzfe7Gb7aRUs3ChvYOMHTFxWQBrWjBSQ
alBF4Jnl5mEVPrfO8ZwqBfUX+PaVTnQLAaJweCRy/8NE3QVKbjzNlw4FTrEY2o/e9e8tcIKVzXpm
1XzredHrEZpeZI6oY7I9OeVEKGFpZbbOj5XXfv8unVrMAXCcDTvZmATgZhN4O7U7XnZlycGg8TwR
u94aHinqpKUCUgwZtfrEolkepHKbVFR9S0KEa7fHaAt+bBhSUFvCyYrN4Kd/ZI1tYcp/lu12ge7Q
WrPZk9zZpHq38hgQbnkbVc+IsvEWUHULsSSIaFua34J4sKlGfHIKjOZ/szpRB1okTY1H1qnGjv/Q
cHHEH7mM2TTWGLU46jN0VXSvOcB2G7qeB4FC5eL0fyO1ezOSgT4L7Ra58rlO3MppKyrGSAGLo6kv
lB801ys8lNcpfwsoo92kiUfhPAU33xJYxL2CZ/nRrunV2KAJlBgf+Eria6OxEhTAbVFzpSmpQV2Z
eYpTG99r6tTCj4J4hArpRcTX6BevS6YGW+h94YeUOUH/1YtoMyLs1uDwzQ77hfHg1dJ0KACANuZM
q/qeK08A4ly34hnDJdu3luwjKezq1FkglJBsFUzGPhj7hWy8Cuw=
`protect end_protected
