-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XtD8ap6pYRPsx8B7KdkaotI7zEWAS8mYcKyT58SAy6L6nL3FenFvYGaBUtgQsiSBPc9csyhyZmpJ
mTbRT5YseL6loj2rRRnEBqLxZb9ulCFAgjR7HKtcMIKeYu2Ssm1JmWS2jDWRNnPLsWJdAVXtR2n0
jJ309VCaC0ZZ+e+fC2N+6LODq8TS29HuR6qs7/V6gPTCJ3rM9QQ+PnMGEPpDU7uvv/JGJty1S0zl
SLxHtH8SDAruNDLm0vNVAmiMnw4iOL93qF7fo2H3DxnRnNQ2IMG/bKZWF/P/htB3Hstp63g5fYeW
m6zSSNg6ScNWQOBQemx3N6hkh0XmvbBymh+9SA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5360)
`protect data_block
Afg6irG00UYG/+5LZ7pJ0WZ0D7UiS7eWV9Vs8KENwUBgr6Da1LKoKyfXiSbyNdj43v1m3U7OmBs9
g6iFw8tCQKbCU05lq7LuvkWLm1ZYQAJQt3Vj50Bmg/EHrlhs3R9rOmx2RXGveRozM6DX5RV15D72
JJ9u5/Bcf+4fEH/bcajILb4JsqnsvilDSZKhv50CKEYUzBWtjM7mPdNWDOKOcoG8RHr48ARn3ncL
mRA7fE+lsdlKd5hNovN69ORERcAvIUw/ZmgEULY2CajntdcbrV92JiNA/P7ImZpseEfmXeiKhW/T
PNit/RqIkWBz+CIqC0+exdQACNEW2Ysxq7g1/K/Qc0lmF0W5p2iAWrMh9H7bphDUU9UDa6XgfPHX
aZ0/a5IvjY4+DyeTQ1w0YTeLXi/v4/5oZWegD9CapRUqIgivLVrVT2XNMzQ/xVhCZjNfnyhYi3zA
EEHS5WP3HOnI5d2s/8OvkKrF6WgPNoSFcrH4j/En974LrcKEVEV/lWsUaHCxTxBs6yxmemO8zR5l
Ty59rgE4B6M8Y3GcWyThax4tvenehOTVUrwxPI8jG70Y7iv0AZ7NxQembxQNre2oK/ZN7FoZKqfl
llwM98pMAPjycZw0o85Y3siOQHYMOhT42DC9m6rRWHxJW2U1pT/kxublXUjaT1YlCIUQLVEOm/u/
5jXImeDGN1t+n4SEXBtwE0br3fYHgchRbYwdVW6EdjyyShdicfYJeRcN3FaQJQuIUYp4do+c8u44
ksspoc3ZYO6FGVyqaSnWsK8hOYVQaKtaeafFhqtv1Zt5AWWI7J1CtWE9112FFs9LyYsvyH0UcOu+
C1rTRtBmXyL0okQ4D4v3vNwt4AT7BJ8BsgSBwyMYwRXSkLR0UeKAATkTMmxHY+Bt0eVltLpTs2k4
N6bGwNpkPXF5gO2hftjorJPAU5TKGBl2s4+r97xSFf1cQOxSxxjj6yO6wJSd/CbcgWrRfDvD/k06
8SOlAkKiy2V8ngugP9a5oR0UqfEivgZ7zCwHJv9TesJxTrzRFw77tRPW80WppM0Gz5G7OWnKX1tK
t3XFg0XfwYWHn7i4G5VAjqTATwfDrSBjbgXcknJlNQh0IjwuahdHNlzC/iWj1ImsJV1NiITngScb
KdoCnSVhWBE1+kVDVqMWp8hsmjdSP99LoIYk8Izc3yd1vVuLNUnteUc2VaO6JmHGD/OBtfFDUq8P
Pl50RMBrQZrzulJZ77qg8NaPEU7aoARkOATzNgr0UngzKm+D32qLYrXQ2slWFZ5KK2l6jXstkqei
DalkhzPVIe7nF+KfhOPnrCnl5bOns9sGxqeY44dmsvl0Gg59Yu8sWVYzOIvDOloZmOB+CcraCub5
gNfP2C5ctXCeOkiRdPROM0UDPq9A2IStWbCpwQHMBTEgWg7+I8ou73CUPCOLUGZXhE3HY8vxeHhP
IN6ntoIqRqiHJgiFVs0jr/UrGR1/pdU5rDSSUm6D/qfqw10E6ZToTJUqtPcEFzvVVh88TIZrIdfe
w7BtjsuOo/cbOdQCJZY35lsPbp6yxO6Ui5NOBd+onqPHBXCm4AZQaOgM+LmguMclqmrB/zM+k2aI
emV6M/UGfhatqK1fLuTS4klF0jOmgAifExSh0XQUnbI4oxrhEY128gJLKa7NvcKrhEKzosZn+k0Z
Q8L867CWvrqFT9G1/dvM3xveG/GPi0SBNs5UFUX/5r8YhFVYs61oDM4E8cVXrL7cgp79Tw74PPQ7
abzvl4kEEHsdKqYGBMUSyxzC5vZJ557bYI612S4IQme+jp8NZ8ZV2iC5148NSktsWEZdChx2vC4Z
jjTFcg4cNZr4a7+wq5PoPcCyfdQ30MdO1i+KH/angkxiB2gfHbdu+qr/HpwHdWLenCI5ReDeOqG9
zLlxJGKAaZmWhZ/d2ewaiTC0jb10PMuAWvypsJEZl3/ewHEg61endKaL8umTPjPEs7sSc8+CXSgc
CmkqVjC6oapDXMTy0qp2Io7OuQcp/W5GsLHz70Jid4sQ4ZJHtp8zG2PmaGmFLtxJJl/NQFgl4cyb
ORcgj3fY7EdNI71zSmpkT5gMn9ETURq44cCwcVI1uGCYyf45dQ6vHcMBJxEd1loUgt/3V8I7EFk8
ejGD6Sme+gatEt4sIk50Wc+boS3cBAinEnXV/FMulPExRDGgOrKGzPuT2saT7pZ1JliN6WA4HFkE
fnw4bkX2HmRvpHi1K+AW15HAizF3fRyjMyE6EoIuZ9IQJOnM9yXlbgAkgaNa4bFIxWNU3+WOG41g
bBMA9OQ9Fso3vQUNqx1R9JRm7jq5TlFYxngKgsVmYZ+GJbQMAJJ8xDQY7rwKuaFm+W0y1gy5HMV2
mBi5epzmbvA67hJwPHvC6XjZzsYYbLYkHs+dSrH9dQDxEBVZHDOrnuYXuXIUb6uvOj+aAwZHmKBq
aIhPwJ8046q62vGtLrKMKXdsY7TpDV6VWYlu8y5vjMBrELbuEPnCwsVgPT0uegnCt3GTFpbujc7m
OFpdkNdVLv8Huc/jpAroFBomT+WXFon1PLb1agwP5tvbbiWY9uFLeIMhdRY2Uw11dB12OEZeEsz9
T7I7s+A8S5389oipBquNNSoToHlxLY/HIYZ4PxYKMmud2TTlnfZwqgTszyZ4BusnFzMWPCSMzG82
jIlBlPUee7P27HmmxNX+xp7SGNFLLr3AFOup0pkLIxucfXxF5lL9zyywV8JZ+oi233r8Ta70h2Tq
8wWTr96VSnIjfs7LO7dkECDQlBTS8rNzYCzRvLVGAp5frzAOBrB3c5M5oBAm17DVe+/ztKyN7YC4
V3co/BU4crb3wLtDHT/NznAXkgnJOHSXKHeBTaHodsAqdyxfP+FFx6I+bs6JBbi9XTn53wkYJ26C
KqaaKVi6rHP44+OjcgJysjQSiEHBVDCLmVv9hD/urEwB5a0OzCr8AbkNyKePYWPmerTAKcXuVxc7
Z/mrxySg6mwNmw59fTtNMqZP0bio+EgAIXqvqMKXN+aXFHRJgPDVYCzXuqd4Izqu8jRFzS/mXvss
S36fPQRXleEncaRJGJ+jDh7O4nve7rmRkSG0ZoKskQlXdL+ovkoQYBPjg0wXgZ0wdPZfrqTo0+H5
Mtv87CijCbaUlf5Q40bXez28TETdLIflmhoPKdW9/sWNw7XWYg8FL4XFHELalQVsDcYVFn5AKsWP
ppbjfLF0Mo07mib8/akq5uepjRiQ+/MLurhOQllI55nsv1tlnLsyauWzEfhAFIPtv75mgNPwaJgq
NM1Ejm4i6v7GuqoSnxStngmNRfz18xzJxan8m7hGdx42q42Ejb7ib+iaBj08RXHk47sSZy0bX1fG
caW9KQvgqtZqoP13drb0O2Ws0+Bx5z4QB9T+Uo4p7SlT0q+yNBBuBL4C68wRixJz4aiW5uPhlvRy
Mkxf7KEXi9nCGzl3RTQTiWpPXdUbRfxt67QBrVmQv2XAUb27QWWaqtqRkvhv64c0y/v61hyO6DLX
ouqpXVne+5ls9pWyjDCe4s9xmRpFEQ19fGMv7idU5192t4N3PaDsOEyMHXn3SH80yBKAoxXa5sPA
tg2Pv2Z1SWRq71JjWldlLtoxsemvUaXJv6rA40KFvPpRj3W4BH8XEsb5qErA7sgCMtdFnwlPE5Me
6w6FjaGE3FQlk5Cx9pz5IwOLuWuMP6Nu9CQwXn87/8TA90Xo+jckMHjjnyooMXxH9SimJX8MFzsc
j23g1lscehGmYVR1j4I3MSPaxf5RoewNows9NwwULjN3v6TlBj+dkoMxtmI/1qlkrWAZZQJ4T7Xj
6gL9xh0xBFKLr1IHoWzhLixVatktRLOjTPn3B/pA+74QkwO6LQjcAKPnQ6GkaIM6OoXBYx4T82p4
mFLtLhKdu68TQKjZptqbbKRtdwmH+EiUN2sS67wWxvxrtsHFAHc4m1g50Mx27orL3tZRJbUGWvlX
mK6HOCimP5Wob7jd39/4Njd5syLpt+OMLxD4g9Cz4PKuapkQXOado1tjsBxJA6vQs2ea/IkKoNdM
k8LoYNM08JsrYR8EHoJBssypjDzvyYQjiBHSAOPanjweZ1Xy4qDCuqFVFmDA/kepMh1pi5g2xKen
uYFj8dM7i3Qw7pBzGAPtoc6P1FX/oUimOiqp2aP4yu24RFm4aBOHGYlofDnSYOe03vFW2bBDuf4V
6A7zBp1obm+wB2+/IVPGQqEee//fwFDjVV/lmVcNHyq5qV7hALNIBNUBHrPFqHmRNO7WykYHLy1M
vEFZLge0wTa+BcJQPJepry/8ju5d5VZBqx3jl8Qq15KxZqW9Y4XyBfe6XSTZ0wIUwB8+KSJCx7mm
wWt4WO79uoF6ChRAcnsGdfss0yYkCMO2vydzE9hzyaSrDEaArPSJ/kdHo9qo3QQpz6ymu7DxP4Ux
0Qu7tyGSAzSzVmfBIwfUnxm/wcT0wqZ9JcTpZDc20/k52B57R42ds5TQwet1EyfquvGxJMvq7nW7
TdzASl9VQ3QnA9dZc9OwvqwwhWpU7wYMbLpAGD+38POsiEFPboJ+KBcGQ2b1pPu0WZthuv1cIINB
zIjkD0JiWcS6yPYp2VmRbjmvfT/aYmuXZirUWNS4MiUixgSw+ehHNoVn/CuXP29jJUnGmZ2tflB2
ZlL7MNZT4RfZBpVlUA2GDSvgK/k6yiVPhXYXP+oXy/uN8XIXEtnvFJhfcpuZyd2LjqWqtGuIScYI
zkmGKxpOaqt6mVF3f2EZzrQJ4FnaQiHn9/J90haGNNbVDUvxEssIR9lRzxF55omMRjcto8rzK4g/
gq5szslC9il27Ml5MSUaS67Ivmn6+94cdSh5Cee5Li7v8QUciTRpNK8QUp85Ip7CYaUL0NkO3StO
BiMU1RfxZS87QkWMsmFZ6UBPEUbMd+1vKg7MXFzq8Wyt+LYULfBmXtdq9wcZHUaHEJlYYMWaBwFt
Ohf8a8ssIZsav/aFhoiTZIL8E1n5oQbZZO0Wydz5+d8Q5w5vddER1Dtvd9Kt9hN2rY1YhLSeFlxs
ofClGSfay2snByMGABd2yjhqBoTqh7IZeP/u9uFtL/Cc+2oxns9z2gkd8XvE7Mb5yx0Diee1DN73
RNFIOuIIGJjFJvXmGLhH+3aIBbUCUvfkLho6fU/LCjBFumv3gxupMOgohjx/izfEXdGAeyjOIkMe
e4QKbXWcvxN9S8BcrOJeUSQrcQGyhczo7Ju/EiuimuHohIGGVrmPgMpqWHFW3rUQ6897DkdTiuAv
IdgaoNcqwzBLUnegVNiGDQ0iuETX+E+32NzEySqij+5sNcQ/4ald8Qk9qYPZhS+2ySNbxiJ6RC38
p/BLXMBEHkDpZyje5zJ2D2zzqKYaX46xOHyyszz+TKC7dBJ3cK0dHb4C7Kyl5w5PAFP9U4x0YeHA
3J0VhcUaEAstXuRNqzfT/jYljVM2s7y79+7LbskOeM3DsZWxJpt+9/6i6Q+ep+qC4B7TIBEmOxNJ
w98HYZnVLZ3BTA2lqiOJ+1RuhoNpLynqY9MQ3OjX5vriJb0z4J1vbNLpnWimpgDbdPLuIt4kSaUE
s5fBCfiGjCeVW5dMh4Q3JS6NVJOCdAP9467otFUKaPNtcZRy90JAH4H1vD6RNXy0D06rN86e2f3p
+yMlilMwbWB/MKQHOPvPHUP8zBMo65JNxmJ4hnZbm9TqF3QQSz0El1ajkBH5O97dD2pfGgxPQ0vi
vg2CEEcf91sclR2WtkI2H6k8J8lI6osH7slycYcd5IjZ3JWiyksMZZ4qaMQsFUAg9uh2nYmWlyvk
wmlziIh8w2H4X4zhxyw8+zPRrnEzr5Xv816EIaob1EiWW+elQtChA/rriQsqOwl8ESNTfI9SuSit
Ifij+cJDGkVruU4ZwlBOzrXzhAqLR8G2QYYn62hOtp6XZiIzv47dSSVkXl8JFWO+CY/urMlf3DCn
oWm2Fz2SrZLKDwVW/VtX0MD7619DuN6ktJkVMT9lX8Y/nQhGjDwLd6ypqZ0DhcXoeWYez3WHZFft
nzh8QCqZnNduKEs63iZMDb18gYo8MscWbcXnRuehvShS/pPq2jupLBW0gdbii+eAY7R/yy0/sNzH
7xVItDX/jkZVlqx09+dmQkb6NnJd/2MZJinYkhxz++ESfdoMK4WWS6/ZqhUPUN0/mxD21adVQ66R
PDeljtYl1hmwLc35qZrvNO5rjZone5O9i4vIOMuN71NwPqz9NkGaR71B7gIIyCHZPnWH90fcS2zX
0TRaWdfWZ4jN5dlBPXBIZbEuJuFlAImLzPn3AHwlnFfwL0wEo5ZVXiG5hFuk1tMuf0YYQLNMbXQ+
OxtZGCWhNAgj0VRPxSxvCm544GQINu93CoPRv+1Oq0FFph4KQeelj6JpWPOx+y+whu5n8/w66kJI
t5Pe9Um7zrXEtOr6YLJLPDP4V1nFrpy8Ki1N3ZPtQT14g0nhzdwqb+900vTfFOhJsM9DQwZgFr/F
gE6egXtCtLftGPkswKCnZPCS+fqXXBIxA4W+VKu4yFFlvZY19L/h60gcFpdZ8GpazNuqGWGsIFB8
1ScMRTYaMFHu2xJ8su+OeIFsAL9dyVUaHu4i5BubqDnwQPHeVdntQVKhNymZs9tkrT3DyUQROHGr
WEr1KIkzv+tkfrfbUt7cYj/hr0EL+KCQfHVviPf3GxKrhgYZPW2kDKcrRubKDCX/lc+2Y7pHnsxK
lA1iYPn4bqK2EeZ5ARVjHxAQsLLftfAMYL+YjkgFjPnE5BkyTKaYkHjjVZ7vNQOIAhxlVG3b8EsT
H+h+RXQio1KTAWT/xORwi7Odje6lYJiswHv6/qyGcwdpuewCv1KOK3LUAuqkPBxB/WzINou3++WZ
PLHvJNLA1bfBXAUQ0E2t4OrOBKEV7wL2UMBPAFe9ZS8t/vbloQboZ0z2D7+2bzoCiaJVH4tcfTaI
2+tY9MfUkvgSMvkPy9mydC+8i69eXDmf3EYQGO+Zal6VM1y2Fx8Vdc+klwMIrcPoO5ji00hXZELR
HG8ZTuFKTL1+8qAtrxFrMhIeJs0+ONdIPm9WpW1vAM0dhBJtpM4BVEVZvk/rQExpiuu1bug5VuyM
cn5ic32CXuHu1eBWveE+10SpaeLKuu5pbyha9vzW63DAdeZjtRbZCgsQfgEcrUJaQDCtZEZLDwpd
j8c=
`protect end_protected
