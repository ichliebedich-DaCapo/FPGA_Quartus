-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lBzyPhqXKhw5TLZPeN4it/b2KOo88RC4UOBW/foAc/2xQ+4j3pjoJEjADMX0ZpNraHMefJrcPJPp
FNZEFCRgitWT+Fbg4VchHYpRBZEeHy3/ei8N0xdqzcbXOyWHkTzpOVSr+RhXquu5WUFSBkQ7WYo4
OkW2+ejJ1T77IE0V+8ks3VVz8wUNyIP5bn6Fv0yy2AQWdMClhwUqmw0PCdBaW8tn4sLYTszy4dPi
eWrVY07//pMIdRRVm9SXSEjS4BfP3ix0ZbqXvxDyzsswWnLiDT+EQjn8r+h7RFpeCAOeldPHUfEn
RzvUlMcAGT9qhXMiKBT/a5x/Ijef2EKquFq0Zg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 43024)
`protect data_block
8Zgv8vndIi9Yy0820cnq2RFNqkCKel5OcC1Fh8ntgOlAznmxGjOBPSKNkr7gL7b+mbbEpZ4fWMuR
NgY8Bd0XTxU6lYtqB0nUSzRRwsnwAsrBQaGzlvKNI315aFtLvQ3sPjbRnJbsB/Kt3+ye2bOBH779
XgZXzBYHro78PKt48rDq0qNblhMM30gcHkfMVZiX7QMawMjNh2YzJ7ZcSIekbJOrhIanbfyLaPZH
MlcSBG0u1UiaKBQCun2dNG/ialdacf2SbyPxsFw3Bnun7pEGyosB0Prydh976Q6Bl65goM+z6OeQ
Zop2JxTJUPocAGXMyv3yjVKiYWxIqmkvht7lkIl2L1OZuNfsHwaDB/I8ePood+Bh3njlqDqxOXC4
QH5XmipwyqL0FInXSWCfu6MAXbYpiBosV32D7R+hJXZDoD7ZEKpXiSaCm+D8RelqTYAuX6ds4CNt
v3qPG7bwyBBLD83TDWLTHzIRexFNIOwBHHjcb3VZQAEeynLocAt0Bjh0H7ZFaEMCr2QWO2zkfRUG
AoJlXDDcgEbNn0xj9OzGLWmglUQUlNr5uQT2e43RXJZoIK1j770pMnDTGfrwPClsBP9k7lzyCZzQ
bm3svLLzM/DE3Llb0djQTcrjAKfYlXxXkLcbLRevRBB/vGJYK7bdpEZvxAvJQn3b/JKmANrRk5XF
1iwgzqhFgTr7pQZ2dtNuLxbgdGpFu/1OAe0j2TgFoyeohNflMsScs5Ac5pBsuz8cdQgcl1CbQnt/
Bef/mOVUaIzqX3nnBdK1VCwlnuQ+knk4y99H3wOzsqhvXBkmGvzXLQx0gQQQg8lLuDIxJZrBGnc3
pU3nwT81yd8DdUHkfWq5P0B43/Xun3xKteMdjEf3F2FWRKT/b+IMv+No4GPB5n8hRC9bEx6h1JPj
h+EJUDAel0+TsWgEndndVsSSbQyiG3CNqP7q+48cmr+ZJrpxZcV2/uvfeoLJmfOgIaUMbogePPIQ
f+SmD+fMCA4Nj5zeGMk9LvHGpZPAV7NNkQXrkGbETogZGw/Bsbkg52UFNjK4iExNmpvgYucfFK7x
o2XCoLwRh1RGWwh3EMzu3O68WcmrSMcwB13rZFsqVt+C27AwLNtXPsNNghB8x8LM/MVbmOBGMX/G
LypzD/wLSpEzMJWzAAeGnSa/73zT3D9zu7wze0lCjEwB+WBVKSSfHmgQCOdkZQ1tP6tVuTFmTZdj
VR81ZaqnyRDzVdkeS1toVWgEav3uMSjbK96igYHbGprE/1xtTs/+COS5ZKkGdWvd66WXpVVM+ZBe
QryA5RLQfDHpYAdjHXcZf5KYfPstirzoEQmt2l1JxHJKRQ+cdTv2chc0J2q9pEfSnX3LqDs2N9f3
QEjsyMs7d2nHpRfhSChQCB/SJZPNeA0CKDrVnB8kWWAxwsIeLZ1GJ9E+iqGpJp0gbebxKkognkng
9p57tnPLk15bKyCFXzEcxLC059HhnFJxnYxqVGJ4HXNi+W4tIjl4KbV8I3dHpB2s/97Hsl5jVvTz
oDbMUqXHnmaoYBkSlU+VbK7w7loSLiV64KbFVZkESKmvBiKPhfzrG1nsSM1PhIMCMitgMLHc+ZeO
xhdLwC29UYcpVwiHSAn1S5e42em4GSJNNZ2Fhkec2uei6BFQgS/gtc2q017Ksvo1PZvzzJpGYx76
DV4GJ7LlMfskP8kWyTGSpQL5FuQhA8hcDvDtNGVRUsa5z2rNBt2rWRFTqSwjeyFTRTBgGPL1/jhf
hyxMLl0dnlnTib5JKFxKMCV09VwORj6xq1EMoceVZp3P8fNTG1e3iGP2OCNoSvjHqcB/28zLOGPj
XHdLsNdn7BVbrmzsPwYSUftTB2ZZqCXPSDlzqF2G9DmR+FT03S+SGyouQyyLl4kLUvzhX592aRCF
snGC3svo31hwIbNfyAMpz7xnGHG033gt7ARIq9rutJM2gzav3Qbr0eSKtWi10HRlIkKIzATc8ijF
7IyyVHjxVV28A8HsvkAzyd0ZYmZQzoW8qsbADnGt72ZjJJeqQlxrHPHTwKplRVZZPW4pACY7j++y
eNspSqu2Nz8draWcvhAVsWxO/UJizHQM/8FDVVNh7vvc9JyHRh30PM3vCQxFzDcvaY5uN5z9XYhN
PZVb/bPed69OINbQ9iCfwcGW9y9e39Ivp3O4ZHCuctxpAdDngFD+wUNgdTxp0T7EurHcccHNl4gs
OS7+OlXv3xG5LyN4HLhZlRkSlSrwRlpwJr1MEBHteTqA5Xg8d+cCwYjD61bcYGYOi+4oAyI8Ifvp
mNJKpDG4Ien/omMEhrqYsv8sxAz7rLNftZ9vJUptgAlCdu0fKL8MvI7Zs9bS4u4azWak4Cua9e3F
n/BAgJBN5Kupbq2ndsSYBhikH4hMj1MmqNNcw7L2Dm3nwvQ01mPbJY4mw+/bnSVFioHurl58wxbL
SwJM0mJa0nT048W1BA5tzbhI9nHd0kAA7bPONnNbvHEoOFn0hws84YlKpXJeO8uQFW2yIcXJxpSP
Yetf/cehIINBKabbUChaROR5ARWME63y52agBDUOVP9Bn6+3f5n9A2GygDGqMejODnkaoz9M0ASs
7S2N4NZpqC5mPbouDaw1dQd6Ep+7i2AY94YDiDAWX9oj51y1imXcklX31UZ33Ji46I3o6KZC3hg9
7JTDmCfYE1UTh7/ISSk59D+zahdv2IGBzGyf+j/YgmQGJh9h9Pne62b/TbZXwIJfPFoIh0N65+6t
vcInQk1nmEGd7vboyrHgDG2jTmf6bJxVSVeMbxL4QJ7hoaNOm2tqg8oqtSi6QHlxQY92ByVV0mZH
SeoxIr1iqJdYcv5ueojFFgt/ss5QN0vVXkDwuYwHuTpTTPd7rVeYqbWzjI6isaxYL5pZ6VvOhWsD
ovzo3FgRIpPnGE6LU6uEGChhsCUxHGo+97e+PxM+8BVJ1z5VsBEC8x/ZdTGD4pVWmWoMMvuMjW3B
4MM+WFiFtR9/rEEmj/UEO81rlNUJZiPQBSr0dXNkOLaR3SYdo6AXPWqPeaAnyWZ9TMw2FhvCR1A4
CMKJU9QVC97N+jRR7AJqBTBZxebV8oXyHQTGkwXRSTmTpSLIXVSoMIROEfgOQkJxMFhgyRUL3s48
7xRccfSr57I3cLS1eD66kbLoH2jrgHj7AlkZFn7owCSFzgbatwoVw9J4uR4hNx6MjozNxnXLnIPE
j22vAZY3ZQjGd9GizoF6cStlRCpV1T7SMJDJnqFE4Jlwr72jvL+81lKv411m09p7oWS8HSNbz7f5
SLjYheg32C55aNRDCqnWaG7zkwRd6BRYgq+4v5DThRPjz2xjgOffiP5px+hqfYY9qsax7EiPN7MR
NEQSBxmwtzKFOKdr8IHFKJ7KPb2AkEEkviod25QqT8xXV7ORdFjZONAkpgS35Rl3+i0WHs+vqsGL
W2EcSzvUtQhSyXsjT/vP8knYqLecJKXUOXpKzUnHzM1XsG09A13j9OTmuzJCorDzqAU68yXXUa8k
pY1WG6aiUitKrQDlENwu5uoHcrQdKdlDtf5pPbjp/jdGEsOUYZgKJb2BaDln2oAjNYMDaLUhyqjM
2Up9tTHQt0pcHjpwhTW2oDCF4pDG4/dDasSXUbdh2st90zr2dCsNtx0mivuYtMtoym6nykOwYVNF
4JDPQ6bUtxilJ2FTktK8hqUfTC9BJ2Qu4LbXVpRlvBU4/VVnuzup7GudHkSFpVNnwJDCzrQsshbk
neDIEDjEau6TQEEpHEz16TpWjW9SmG8Ivo/yLko03jZ41RIJL6InSFiBUURTNbmoSCclo8hW60FL
joIKN0mcfOtTarKVdLsg+lFpdHcADrvPtlF+/9iifZWN+m498i0ZfLcWkei46q6eePTgMksE70YX
UMu+gZx7hpeSiY3bw192GbU4DbcdfzXNoKiJbCrUD9jVV+lHFVd94yji2Qk3FNr5sYmOnpBIGbWW
HZLVJD+3UxNKWv3nXV8QUONygBCWuPO0mOXJAHeC3yDX1R4rSsGNIkQyCCOKDbvQBHSiT1ZTuHC8
grVkqTWxaMyoglHd9bSG0zZj+E6287BOu5PrHxDIqzGwdkAyU4Hfv9s+V/T5V9PiCPvm3b+aL8UR
AJ2H8eN3O9BrsXX8m/jqr40Uz+wQYEbsp8bqQ5CUocnzBG9qdfVQZEkVuMiC3Tgm86LdSM4YA6nQ
YIl2IuEaKNvbhXgpiZ5Uzpx2BoJ84Bi+CiflseqRLcUGNbAysgLXoIslltOWnJtFhpFQbPPHIk+V
sb7Gad+NbOrK2jz6beWnmkOB2FzQuyEPUNrlyOYo/e/JOdjLf/tF65OOPy7bV3A7voOery8OkptA
TbnLRjuvKjbTlzwtWwhk3iNGXh7Sm2LjGKPHLvAHatdEFx8n37sEyHEZY3oMlMfLvaD+VVebnvNL
M2Eg+f4cy5lU/YCUc++l4YN8hfM27khY5HRvo2DvCDABb69/bZdPbVOTSHdAoQs8tsAH8/ydMvvk
6gjf4PXOrTGt+zcftr8wL5PREgSv7/aSFmY7VQzbNN3q/RJ+Gd2HZw4lMzhshbt+w31bWYoMuHBK
3soe8GFGA1LwCjyrMZtE+EA7RLSkYbum0zOKoUgr5S3j4wnMCX+FzjIDjTtWnyycR9m5F356lYDG
cGOYyjZnqmhH87ZWPCPvfadNmMW061T5sjoFgT/GeigA8IbO0f6SEMxL6GpFY18EMDk33Ke/eTJu
AUiOM/RI7dUUz3E5vyx8QUi/ddWmZSoMMxJLxCQKyEkwHBmyjcKO5JE+OZuXggJKNjKSsyMy9Gav
BPuj2uxhbknPEVWy0frkBleWjo0Cz+tqcyoSLH/uvQTtQcStgL4ylj2bR6nfUdjzukewPJr6gkxM
0sF1kb9nu5bk3oN8vS1CKp8lBCt/SSUdDmJIoEr8WrLXnJRz0t6NsyYxdRTv2Yat6OE49NPMGecs
1bgEaihnjfUSZlw92xdZvfHsVBE9lE62W0PgGpfnP4txsML0chr0ooojr4uq0VmQEjy50tWN9d8c
2JEfKLz/f2XieUf/Lg2sL1peiw6zhH00/6EhUnSUmpLw4CySS1cVMPcyWDCtTSL1nkQAvWSBuZPl
agpwAgbgrmO1OO5KxPGvToEaKwza7EN8yvazNfkDxY0nJH2Lg0V48XHDU8qG1XmIU3ss9zxCSssm
MmSvYtRvul4bG97spyl1fwgEMjuU9SbZ3YvOX4mAj/6Chg3vRVGfzJpzbG98OeOtu5W39h4W5qS9
PqNkI81JEuoaAJGOhDSFaJj3AdkE3ePu0FdMOmgznoFIq2tsLzMz7EFBksy/ZA+iivbg6jtsxsit
PfW8HTuVgljAFjUbqR2wWSD8tzJkTm0r9hHMzjEBvTeB8z6d/3uxBt6Qluyno7TkK+gjosHcJKHw
X+P+eik5Z6Qg55pBz8g+VssoxW7iaYHgpUsR9geOyqarhuZ8Zz3hBE43CgLXP+t2ogMCaBqceWIe
WAZiF6/xUFtxY3KBNhvsrluJaI1LPaS8QbvgFx6esGYUbF3gk0KdOrQ+jDBA8vl4saYeihxDWUzG
1HOPP+4mTiIqDGe3tLtJWeN2OvmMzaKz/rlMBU+niqhrHCHGrKr+XW1zQcxoPe6o/JwBUOOgYGIJ
hQNA8ggG/bINgWIO6UnCKosXgRdCdYzS6TWI8gaO7XR8nLzqM/gbiRfoBrN/6uPOdA67hdKqnay/
WgdZPGUaXG42TcYP1Wob/96yS5hZkPILSr1JU9HSoAKOxLyY2PXFUrA84V4JCkGuwr+vdVRWtOeP
Xf0B2jtrtXKdvWsEh6FvTevfkcTXVXf6Ziju0Xpewv2MRedE5IZXPvUIz+CEkX8KTCMAawCuZ5Vq
xelRaYDQTDV0MDkhSw2tAg3zp5IrpbTdD7kwOiEastGMTZMCT2/myJhJZfCUTUW2HP08z4EZm1be
rlAcYHPUlA3WsmZpulU4TwhrsagRgXwRUASlD6LZ3I5hYHZbttw6F8v7c0qX1qiKLhF36wAUlZCX
SgiMcJ+/AvPNlbHl0xJV4JdyuuXyPOBkU7glInbMViWrXkfNnWFIJHaOMNju5sa3eOlLXj/eASrs
5vI3REp2OMjjpS1JqDQpok9JamOqGtKb1RHeWPa9L2AcgJ3yR0pBjVIchnHFuzgcBB97elt93LRw
26lIU1UgSTQdLvDKmVTk2SVowLOHR8BtOombL5tTfIrfyod2mFOVJFbaAQ8VxHfh1Eozvh7Z8bm/
CKss8kPoBmCuCto+jHuL1dnKUiFBKH5qfVtbE5Z2L28tdK2dNUpsBg6XL/vX4LsXj3ve8P++LrCl
Khf18auJ8US/OGsn8RqGg1uJDPg6fvoYBuUCrKyPGLPDZhXgJtpuWBg027gkH7krHoKORyNJZ+3h
LOo3+PFsOCaMUk1qbjs+u+Nhr27t8ig56h2pQ2ho/Fiw9wQAy4Ilr6LUjInV19rgjKBDOwvc3jmU
/W9iQGLzFG4U+VYHggpYwepA0SMr7eFq46iTQ2oIXoZqvsMZ8u4WIKJbUyHtXCajp5SXDKH7ByDI
bSWYfBY/D1x/bbz4BWIUMYfU2ul8qARJpM+KMR0X052oVXvBfG5kccjXPzymdYGcl9bvT9/OYXMZ
fdCBVL0JGvlNdLZkzPGJ5IEf1tg+Q1fxMAibjcQVbNQyBSnwgZo9fvjBrQRPESUCEpzB99wH9YUC
0oWVPfxMjt5YDbU6FCo6MkPIFSPknJn2mE5lnhxsS+wex2ECtMyMQKgOtcrIqFLsd5nGr7D1bYp8
RzIWXEje71WVmtgWMgRrcyiKWvy6dnsRVZB9IX9xma2PUqBPhbDaqmOg4UYRsHKKlAEA5CnU9fk/
aKihlw0vRnoN5Zqa48QEt5bhmnPrzteFPwVchb7YmkFDxekxE9UDjGMNC4Av/wvmo8lQG4Z7Nihp
ocgZC7ojd7pq6Um3A36sz4m+icwG0bitiCguvlpvBe+aGFsSxAaahTFgAGU+jiWVe7/i8kGosCKC
MCQbNphUxvJOR723M3MaFYgaXq2gc0OTJQ1S9rFxzzw8qPbzLlIsMDP4TkMA3cqh14FRxgfxPPuu
NgWilJe270QD19j3Z1lD0nSSqriJMtFuqKZE5PYP5K6g0D422OaKcKGB1PyKGyONMZ5Li7sylL/F
bYwt0uZE3H+fGUe6wm8idSmfea7lo2IkELxHJO1YjBKDdVkELxt0KsAzP9jkOiaLo6ML6H2Yv8n2
nxLA5GeP3S3bWg3VQ3FezcyQ0ccgIRQFYIsYHooPrvGcb/oJh8tyXf0CmdwA9oZM/BMPvokr4lHJ
y+8yhjZAugq2ZlUjiZDF0082vME8/qyp/IR6HyP1LDttX+tWW8WoEuPBz3YbgE52GuIrTDcxxWeb
TTb/kmo8b1yChKVPzh74k+AL2gDLi+OOXEtfgAVXtbnboxs+low4v+H7YvwkLMgWU1rhMWQx/Qao
5jNkbHwd/fdGAK883itBZVrV8rkvninrhc/OXjPR/6v9ULnSOSFggG5OXtasU5MMWOgCCcXHKx8p
IZJdZfHCCSoSxgUu2GejcnsOxZUjFdBlC8/GOpW1T0idG+bfonGGmzgj3DEAcUWwkNKgqurqeajb
f7/iwrGvL5qXKgcfj64NjZixl2hwrTRoOi1/lI51RZuGGL/6CeJZm6fhGMU3jfbaWBPseyUj2kVk
ng7dlABS/9A10Q7MQsY8MD0AHk1I01XBp1bkBOi79vSRDA2i33EYqGWvgPbQKtvMg09p8pfxwACV
8YUyQJEvAH1pMdvv06VusvouvnIhg80x1KxRMjL8MGCkP744TbtG4ocLZIjP3N3i9LdZ/ZQxC9UV
dbNTI7n+Tq2jhMeBl3kWrA+pw4EDA9AE3vPKF/RvApY1ScQ507dUUBZgiAULzR98RLCP3EQ/TmVU
MGTnMzLwy+HJ6MOLny67uNSSgii8ZwC9fqryitjLmXi1m0C8lNCfHeQm64fbF/cpswn/IW0szivd
5alJM95UEl6TNsbaeW6CFqQSjdHjdIT9eGB6cmSIzhhktS9nhOooCaY24HuWKPwuO4o2J+Y8sgPN
eh+oSov7qZ7RJADu3LRvXYhBrBbYrEHc//rgxzi60cvxLz4PxmBbZbYEJk6CMyZCKrSbvRbpUiaO
qb7rmIvo98VL4CrOs1GYe9QrINl66+fvG2aY6TnXBHdUMofEsGrACjKBmMkqrxUjMX7KR8Br1Zvw
t8WrX0z38pvjHWkteH+nEPcNoPJ/WRSlpIgeBTU4h1hAKf7G2XtbMcDnEGLQSN9qcQm0vBG27Toq
OdNN2tQXE9t4PViiKTH8+zVBWKGOv+/Qm2Gu1B0wd9fllcxHSkIdmHrDd0wVIZT+AGteP+Pt6wBb
coO8d8iSBvmsnhzbKqxF8NVmhIeA6E76iacWTsXIKfDNRG74eJ70+/HKk0zNWViCjS1SLYQJ5KMW
E1JdZS7ftPIp5P+R9gESrtIf7H8wt/pBq5lFrCJZlZgAfbZEtIXtzaqfyzeSHwE6KFuDdIasqvDf
L96/Hr60bsp2iIlb0K+60a11YPj44xeYIAFbvVoQ2GQXSOI/g7KNQmLR3YXxlWRBvvqFIl4jX7Zw
sRE9ZL/mSzsLedSISUV2W9ZPO/+N5Q2ZfHITslUKOWJKa3UN2Z9na4aKMfWRregR3CBPkP69G/5O
ceSVTFVNU/JS9nZ58evvtaPahBzYy70Qhml/NJRxC+zWIASYs3eKvTKxi2m2nAXe/iV4GBWqWkdf
gQg7P6VXwKIWzYXQqpYy8mxZZr6FZZPIYxSob7tLtUqVU4hT8PrKRZcrncNORbvJgqMX3Pno9oyT
pQdcYEt2cAepCWttYU2krklQeKYlc+xZZNAOLQRN5QSHrPlxaB916+tbU/1y8X400xeXei6rkvUa
b7UPilsxZLTUZ268umaZ0zrPVEVn1/3s6ovgwM3s9jhoRRH9JC7hSawVMHoLNRkgvOoAs71KLVH5
x+6xtxtY4JdSA8uIataefOvlDDykWTYs9ZWN+qSz7QwUZ52Gheg+koA6rL28DWiB8NIFb4GwynH1
UF6hxzVsvV02TuQDyTG/iu7GYjehuaP4C5WF5Yq6QNNgl+n2VM5a5al1IDKMHCHH6Lpwaa2Nk8k0
uKG1uo6hYeqiZ/mg5bTfBzU9K20EGxxLxacyRrf/hJUWHjFlJKi7QgFOVntkjjtMVvDAAqvkGYLA
qc10J+0TOawvn6dXs4fr85ARQoPwS5kxoZxrBWvBLzfVVO2FZfapjBdxZjTwTt1ebRMegCETYfyO
FmfWr7S7shRP66kxTFhKHcAkzGQmP6+Xokb/LDD/jbI4dIEa9ZilBThaf07CvsgORYjHA6l6Sx+R
F1yKPM/y81zHZ2w13nm5b6S9QqCxLqbld/KVLEo/wfMykUc2CCvb0OBCElYoTyghXP3YGqqZemNl
q3JnK0X59wlth6wGieRAuvEzY9OkSWbPnexJRiLF51yn/vB12LpZ2CuNtsdqI3coN0e6LfUFmx9Z
SAL1C94k0SV+TFkUn6c9vAOKgmTGZl987oc+fnwCUIncaqewwylLQFgvAySStUWR5lJz3sUiPPAs
5UzfpWwnP6NETIx2hBw0sAw/jPPj59PNMEDKGu5L3SPacyqrqO1e3ZIeceKM9c5dDlcduubZkwaV
mUWefcES+N+mty95gQioHI+HuS0C6sE1O09G4Cv8+ayphkkn7/knoy4oCuYQ/eVrKyQsIf+LMSf6
YjJsc8b+7LdXvzg8+ZrnWbHMhKDCJNFMqZ9Wk94zr8BqDBOCb2yC9A/DxEDtpVH7/WDrGxa/X3KC
c9QbTwN1ROcJtyfC5gTkmMoByxaop5XOiFsV4aYrBKZS2bfpaa+5Tfuoo6EMdPZcsV+7psajliCQ
pdVIzlEUFNjyLhEpX7SqqEaG7HjyCYv6HItiB6+o68ZibK5WgzatQKJXAeoGzzE1qRfJceCtCg/U
aveRcG9nx4st7zfPUuh9LpQMhe0rNXziy38BLZiF2Lvsxc85zYxk5DG2ymIh10+oJTWDFoO92CpL
LfJwPyDznSSQz9M6entup9FqMKGrVxw5JPr/8k43Acgseror6YAWnJuxCMkGXf+Vk1W3jWgM8aVL
Ao5AqIE59bKCJLu9ADAUsbB3Bh/KuDEPHCBeHiXsuGm1NHTYic+PLnuy4RoFJskeYj8mxUauHlIe
Zyo4TssxdD4s/uSLH9clMXmrwdxUP31yjom0jMmn+oHd2/HDlW9bCX/K2UE0Iqe5vE90t1EakjEM
C1sPaQskf5fzwnNd0g/31kqD+ALQLW/NjZ4FfAJS6BTDJQvraDrdUnJDAeJCQ76VcWubQtOKQxSQ
/Dbh3cOZIZk9xJdAXpfNU7hyKruroPldl4IY8JUYquik0BdclUVyqoPtV2Q2WvpI871R1nmNoXfB
lG2BTHhEyyGS5bN2AdesXz84UWLCVylPOn/TZ2ESEBQPozlLSbdDPatzZroEa3KP0DIcmyfCHWOC
ALXsxmfw1fE0+W4KqfDpef9osBzLqXGJeXt0sEHmIYVgMgH66OWzx8JbcbgW1zjer2Q2idz7GkZG
D4dgfzo8M5L1q6ben5uKoXIY76zkAHieIUrGR8ng/ro0CxHomqhDUAwTP5yXgY0Meeld8ndSEN9z
A3kl5+e/DEh6lr9Ba8PA4eqq3LdPPE7lbulbiIBKIgmA6uU7bw12yOrBdqqsw/Qhs0yBfkXylApz
VkYm5Cdbpo48aN33E5RXHZ7BczLGsVbjWZxo5A3JVAbmjEOpdc3GKVqkAUYW8mTc9dUo9cwZ5rn/
7Idc6EKqqnClp2wQHmCE6OJInzCRAFRuwHHlOyLh4wXnyyWI2jk1aEugn9kAoYegSOwNEuKgsHKp
AsnnzIm+Mih0ds4cFhWy3XEyYHjXNIeQwH3O6MODygTPdignNEm4sVEFvx2KZNWgvl/oaXtP7xzc
g3ZHDpWm5g3SJcPUk+Nww5OXu1rf/C6gul+ASXQ2zjko5LFEkrpaINmm3RSxGOvFhwXKQZBphXbu
OCALMZi8e+NFJABG4Ec1ltJ8uIrlDcv0QMl7cHyEl0ZqMG5Dj1TCtsc+/dugnjDien3RaTTAmxSv
OUC15jtFS2ZxtdqE/n96n+04N3WahJ3MoYljXGAnBs0yzhDdVKQeaxgYO1oacUmqL/qvL7zR1t1L
nrhfaotQS7tS1CPV5hvdXWdsGO8/zJhWnQvwELou3pS3nK5AusnScMx6JqQ3pT45H90P7YKkKVQ5
DJDiXy5l/d1TaxkrCVnoYHd3rTBNGU7ZA/5EQ4Xr4P1QeODKed5QCOCxQFtjSvywS2cqaJ0z6cUh
m/KOMa/BZcT6dugiHhgrseKip6Vhw5N950Kd0f2CvH/NHEUVvS9da6Ip30zrtoTe/2agbhkF8+FF
u2uSwaRO9W2jgfT0ABriWhTcCWaXOlgPfks8WWctwnb6S51LvbxBWLkmBkEJw5ZycPiCzw5r372z
UQSy+dz3zGD89/bw0K3Pys8bADdzltXdYtQlNROLhXBFCrYFFTexJrefqll3tvg3MCg4v8A+HP54
BFy2CZC+TtDivH7zFBHc5x/Hz4sNDoT/NWG6aD57GaoLcUKtMI5oHv/smm+cHIZ20U8CqyPwgE77
DDbS0ISyI10XwkTukRTpne1lS7RU+1nXHJ1h+PXGMUlRbMk2Uu1PsbomIc4VrIP8ID8pWZ1HWhH2
XJC7FU2NljQJbrs8+gOxQzmvPdXt8jDtkbLx24ZdBIz7swOp2AeigB0mEEPgltnO/VTbgcxXoM7O
05fsxqDjjupIfvVdfL9+Cz66nTOrtSBduZLM1DpR8iQkMwk46DXRSJJ5o/NvR+o1yFxfdEsAxUhn
i8szBCYUB3gA4h/4uexqX9XBpPWJIsMH83/IqMPm45ZGEwX0q1t/Lfh5ycG+quRpr6VZ8csrF6xI
J8dvkqtQgo/vhe0l3eVV0fbZkzaKybrJxqzmJKwef7tc6EkaDadHsnOW7cXnKed1K3XWk/IqlK4b
O0MJnECkL7et/5W7mOUaLcAYO8GOL2wdiTzJ4ISwtCztVd1FqFf01UEp8b+2RUndt9548yDUvWRb
YqSx4GOwqmhVQ8hckUaQz+YYEWmGIqjnNPyQ4u9IRPTi/VPd3c844OT2E8RcX8KDloAQfZs2YwKm
qY6wRAeDtbBTESP/Kd4McntMIKo7RqcTOS44sA2rwvj66Ns+HjfxVfOAipLwklgkzsdk1KRcpDVO
PPO32rYbkDJyUfwQ85SMhyU2W2TY8Vmq8CLuEN12ah/SVZoa7Gg+wPjsk182IKlYNYatAqijk2rC
CgmTFwVosMXb81TuX4V1zfs8oVuaMFx8NncIh2PrfGZ2ZbktF8yeTciTaAGk+dRFH1W2xI9ZAG76
OQV3tgyTlxXHBKmThv4Gb3PshCIZgtcoGTrqHIe16eeLTSZ+jYambKMx7wryNS4IRzRuPm2o0XFq
txYPtUySqZDnDFbf3LWwQLuHv36eNMKIZ5GxtFFLFUieig0sxoaINFxMROmn4O0jlZ8ff45uRZwR
hGxJL4D/EGVokC+x0H5vuAnxzGYwNhQvBZ9N+wUWWPYHJZRmNzgsrplcajyiNZfUVX6HvgDIP7Er
/k9YioCa6ZWRHdR9Z1TBKgQ9FLAVt5Poj0zNOOp6NT3v4KxGMXIYlpOfytvfgDblazw0W3BX133+
WlZ8xpF4VwLx1hww2nSHqyiNwxIziQ25Srom+M7aF2epyRXX2nzcerXqJ6ANarqZSVX98Uaxpoi2
h3igfUTfTZ11pkV0h2LzXcUz6qin04XKq/+YXtmURDuWVD1odaesB70Ta9OwVEPxoH2heA7B6Gqf
Ph0v+c6HHtANL/f38Ob+UL31jbp4zKt3g6rLub/yycVun1rr4WfU4lZLHtQfSITNndHYaZtY6yV9
aBqaruNysLK2klbpFbJgNle9kuxWOMLEv9DI+wdEMAtwlI2MEWMqRBF5hABnGwfwkKdeA+X+6Iic
67ZpIN8FHG/JHPYNI9wp5y7gBaoG2VWnUORd/802d7XrUX4a6bk9bXwfBZ5kl1BtAZu5bymZW/k0
jyr3gE+c0bHdMh6WChVjd/pO4JnfKLzf9POtnOlsoHbXv6Y2pslMRn+9rRJm7h4gXpRrtLrRSZZ0
XY1m10lVKpXFEy4db2m2mvKNO3EfNSIlm4U7f1OP58vMyiIc/rKsg6l3dpfxAggSRxokQW83JAmQ
zwX8YSWEp94gQ0T19epTwl6PLDZ/HL60kk1H48IwOf30Kj3ZbiQY4n4VMw7UOD5NzcRSOFD8XwUS
i25MTooVU9l7bcS52APSNHP+NCCpFHbE/+eJFVpV6fivGwamhWEn0MHrtVWvlFD51RcUThbA4s+9
JUGqpFuquMXrZggu/DfAvt+joIgoPDdgpeH9KMMdIJhTLFzp5Bchqi6xwD0rEGUEgd5LYPXVFzdS
N0lOTZLimgEFXu4wT6FMxVBN81OwO4f/5/0GDbaOXxQgLbrAr8r2Of/xK4/m0H0NF9qjs9YKjzh4
+nfe3o+lgymjJLfffrkU3LT2DjWOKxWLd6LbsFvfOgwgphhBuLrnMogfn6//kcpZ1/T5bHBAt6HX
aHj1Vw0CFxk1cwy/l1LQu+JCPUDG3+ksVuHZVhi32kSEJ4oJnRvUE3Yimdk/FZTnWFwbJUnCXYt9
8cbY3jRfrk+4zwk75hIUEcuLprpZmSIfVnY0HMK3R8CR6ICDMaNVf3BGdL8fqP9u2eG+q8eSlcCx
L6D/W1HTGTYBHxCbcgqPn/CsiC6d3LLWi07fewdbuEVax2etN8xDCw7Ka5d0jedQHytu1slCTAyI
EVtG4Yjy5cTEdatwnXT/MjFIPi8Esmt6EpiIejosrM7y662dJas8ggbgkAwbQsJnoiZOgMjvT87Y
oTVgxzCBTnmXCnFG/VWyVMuIKL5LzTREgZFf7Uf8eDIkQ8Cn0GbyG3DOnAXJhc8BABLWNgj1HfOk
TzIehs0DxKfrjJUCTmJ9VDiTCC3IESkOW7+CbCAuEWgsOf5ISvgN2ItzqDa+ALNrUCuTh6b6qtIO
OXq41qhCfGLdAjoAGlIWw1K1iiYhJJ6ec8EMtEJLuLDUp4cUdVtS6aSSwOgw9lyLnFoEbtaIQp27
0SNgNfFrlA9fMmeEFJ9I5l7rEqsS22z2z9oqM+kzhn2houZcTHZyYZMEPno0URaf1fJ3XQNucjM4
oqPphAVH/V8jcy4HgFVBEt4CVAAsyVsX1Ub7gxM+/rgz4TbFoCfKpt4xCf+TQ3BAap7/eIBR8Gdl
AGDhG9rDcl7r0ShPjGYlDcv0BSA4XUTwL+mHWAhDRoOwL+/HeIjm2fnkPz3lr2kaT7GZ1mYlxm6q
r9ddkOWHeHmUV0gaX3AzW6ezvGLruX5IQKCQcmtc65GiYmHhvhXoYi2DNz0vJhaVMSCdox5KX6CN
DcO98inZPbbRSKmkLcZFyow2bt9CIr+5nobIRt5uF0si5uNOM4stk05a8ZV9ACDnplMQQdg6HG0O
OnW/ZF1xKXhneN3II+lbqFKuM9IlRkh1qrfmg5yciIvY4FKFYSFLN06l61X08bDsOEGOsWKWFnbm
pWbw14jMKyoho0srbzCOFT73sasz7Ikl9Lme9ZFRTpVugYnMuRlusqW1Ihc/xxMzzCSzRJqAJY0H
PUQTkP4DwuJR2r4UPAcDir+8Hlh6zofrRhgPExWSz26nmkel/cpfPoo0Z6FNQBRl1akIpP2KECKH
kVMnpvx52LCE0dK2KIn+TYl9LnelJlxuUDXTHfJWJrjBUB9Wl8lcP/4e+bs1NaMQmDqBDP20MsTD
NkQqEGP2n+SG5vPU1sXM027y73gEtmGbKYbkmLy/DuvDi5meIetv17D+LExvPLPp9d7UVxUJUM4e
dZAfXeVPMTEXHpAODNcBw7VwKBWbb97sp0ny/b3Cx4pP7/3u8NOKXEzr4Y7gShpC41l5TgSC2uk0
D/hTVmH3U+0ZGEw6vwftfOVsyBdY1R8aHy0uwpROfuLfXXYH4I01xKo+z2Dq7UF3wroYDh6BPQ4q
1qPBGWBFYD16ympFPC+H02b5QlJnZaH4whGxpZ7ysrBgHEk2dNhfPRvFvyPXRJkyFamvUjVKzOT9
4ABv7Ty1l9LCpIaNwpyoTEdzn69RixgUE/hpGx1xGJJ0BZMJcotQQNizUVZIymYyKyTIs92Zw0K5
4cE+vYEFRGvl4RA1M/phAnv0XqBqJ73StpR/NDt3F9iToNWaov5Cg32mlT0HFdg3pvmllzQhLuXg
wdHIMR+/XoO3OrHCQGbN5cf4mbxF0FH/jzBRLq/yTUk7IAx8YBtL5yfNrnA72b/GFGnZ436NT1tR
vWhGXAJIxGdYNHVGTMIIKbHwxeVIZA/8trgVuyKTngUnlDeOZVHUeo7D9z2krWgfW0fX459ftRIt
TtDQ/iz92erMQ+ew+axhJKx1gH9vHhjV70ods66wggAMdBihAwf7nosEUS/KNFIh3q1wp6WeU7Le
c3ADxlv2dWcZbP+3J5l4cPKw9jDpLjj3qjJXYS1ji4PRylp/8Ij5HDkar21ygsbJOSVH0C9ngbwV
pmCp+P68TPyJ/Ah1IItDrIdCWCWfHBqXCykJf1Hy++oXfO4ShhToswH+FFS8zGvjFDLulqFJ3TPL
ouTNidAFRDkz8mnH9rDGBZka7VeKMu9bgEjlw/L29qJh/0XOjYt12BGu+xannRGGk2svyFp6owZQ
n7oYgp5DlQwm+UKoBawUCbevR5yeHZYW20L24kRbG5N1dvWGrX90GGAyED30i0lvx7UTyJPP6PAw
yV/DJwGU2a4GuLa/uTe5s9uRP2ZYhDb8BqKwz2b6jgXssV0R4vlsbP/qzbGGOoJa72LbZxm/r97z
WnUIFUJOW1Q28Aa5zG/iicGYIOaNDy5MjP5gu4lqn5qr1lKf4AGPjK6g9AnhIrY+SfrUGpj/ubmQ
Tq3MRDkuH6HtJbDOQmFoNisBnvglE2aqZXccT8ufRkvj+38JUszzgHCu1aD9ALcINccOhsMW/XHr
B1WBmVehrUiZj0mpJpQY91/suu0AHplro0fBP9+48wSs3dVnZGZ5lQEsZpd6ZS+Nutj10nU4UuvO
ZDsOafc3TjcK8/Qmdq0k7PM+PxJqyaNm5NxYtkrE9leyyk2MAeqiZ6uiMVI/NgcgWzTlfrGCddWm
82ziaSgLilzQBm0on7V9KozbyUmnLXP7rNfJFin9S+CHkt2Xz/08AoWoQCkScN7cuPUBjqUmJWP8
ZakEMiVdjTd3KNH8ydrwvQeP2U3b5UEpVuY86wn5O/4ZnGtkVb44nbUIu6OpuI8IqXssaVxsrYgy
fimtegjHnylGsn3V74E5BYOpO5TLwE5ykSKTB4gs+HsCcedI7hUlOyKXJ3oq7syQFrcHNNaAuAwH
fG5ntCT9DMRQlaEem66M9DdGV3i8R4nLk6uABuQZQ1bUmuntJs56LqZrS24ozJ0LVDDDOz68jb2H
AmB47HRiR2btMAfNtfFcLGIrpla+n0zxt9X1ZtuVmCYby1thSBPooHmMInYlaeNEzOvLKfMxJsW+
hA7WddPGkzQxNsPfxtWT/WhRfuvU6iWwmiJKAz5Udf9tfBpUOyOBdCW7JAD7DaCuKXcCr4f8ABMD
tgyItHhESsRcmL9pSH2z8XCIwSM3T0pZqOS5R5y0fQgUqJPv611OmZZMgPcnXh7dkmfAtq9izVG2
nbBvC/Zo7zp+X+NKqxmj/GhaGgTdHv694K3A+AjMZCuxbfTtLlgaZNmJqI4F+aVKMkdMIW9TTGJU
Mu3nNdhmlas8euaIb2qgmtClPLZMBgFZUPIrMjUTXR+7vxnwbl2sdgwchG0EkaOSYMrpHstgqEMc
BLVuzRy6xJfTMsOA+Y+QwdhH/MAJ6LdcFIdJF6pOgbfLMw2uQ2HKX8PX7l2VgA6vpEERpZq2Tji/
7NiCEgVOtKJakK4AN+JHqyO7GCeSARimlHZNHyxtUPLeEMXFtyjcfZCaSE/FmtDufkjeCTHOEPM0
gn45PDVirifYeebyfAfe6jsxdLQNtNkl85tQyAEIEza0Skhy+i3f039Hi88XFoOc/Kh4M3wcQmqS
W0JygYHhqtHy4btTg1r6ZR2kA28bZY2Zq+P+d39Dif7TyZtu/eyiJShkpEQeZFjtu3W8JORuUdDo
qSkkS6BQPhBiFqi3sP9R6EXPbVPWMOROUT+TU4uqLsckasZEk+YfZ387SDSaNVy5tgPNGyb9jOD+
GZTc7b6NXBrwwdo26eexyDwKITTcUwhzgNIm1ocKFJ9zRo7lN6V0UZJsLCBP8W5RIBimqGY65HRC
qsdUa2wfYnhC5IPinpcjjjfFarV9F6Nz1J1QnR6EM9NyC2NilCeTr9DlTDzaRe1RiIyKxGPLSlIF
abwbgr9mUaM/+ot+NBcXYsjqKornFgXgfs0aM5yjSeDVUAzm6NfRhD7xbzMFarleHxgMixtbl+U4
uzcul80ntuO7b3bHP+br+TobaCL+7d+q54fKRU2xw9Z2nrrwSJDMtCN3f0gDhtoH9Ts8UetinFao
KIUwElfluw2PkwZ7NfG9sNpkA7VSsZGpacnq9vq512rLDo2/wbsy/+BQH8zsHe8w/zfJxd5WZ3tn
ZdFNvQSAwTYqhNh24D4+FjxpNsGvxGO3YLWAkvKWRABpdRio0TQH5mHLqiOjo+1vcuowIbRPGsRW
MA7A39ySN8aypOWt7kJhXvjrufahcD0R7SXtmaxZM1uPX0PguHzxdu3WPwj3ef365CU1a/tLTEu2
ultrvJc46ic2Mis4QlRB4x0qNVqXEh2brkj5+t+T/azOlAnNrxjtMwrjuWBwojk3rLlgvaBhZ4Fc
PxjNIZtATNK8etGRaoViQ9mbRLgzHFUeCQVg63YJF8017rW3d53ufpyHxUvVdE/NWwzNpmJsLFyg
lm4wnBjfN3dNJC4a7bMAeMcBPcLNloZFFOCm7z7ZMsech9h23dlOqj0YA4CSCWNQvtwrJSXDg+XU
zORSG8fVGLs6XS0OTAPufUPqTOfQORLH1DDS6+/hNEIA18keuL1SW+8Wn6DYcpTEAyPCsUglbqoE
6EYcQTFsPQDpTR7yTFHi3lperVXRCye3wnzvhUDPYICwBaMh/1CV8MBQMN9HEve5wcUYkrsihmlK
hOPl/lKeGTqngXA1AbMT8eFlRTqtARQ45+r9sprShqFSI/bue+NILwOqxGOUF+cmskRL1jS6iXN8
DlCnLgesmiRmd0lrp2chqLEgbwpTwwbWtdVqXGZyA2SMZr1q2PcESzSLrPvzAmTvLF3fbm1RW/Sq
od8g8EkmN6tT3RKMfASlefm4AlT6lAU75pTEjvuji2hHoAOIrMSHi91XOeQ1nLSNPBD+Ck0qkGip
YUQs0WRWvrc503yc4tTpO3CGQRIqxT/c84tWAgU74zk20uYFs/JX+bSUacm0ba8yY49Dbj9r6myk
uSXLffP/mFgTdAFz+bj/0DWveEkx6A20xHPLrsDGksKFxhsGzAO5DfOvaUuFxV/YqallaqOxxJd8
deGk4Cy0OQRGQ5IYKWWkZXe6wRFrpUtvSoqkaGxephsgCuJP5DptecuYohiAXbOxG+MuN6mE+Zh0
PzzBclQNFcNDhwtIJMiCW8o8/tAxKs8F4woapJmg457lCZxAQfkSYp1Nk4CDLC38NyWhunaSVOX2
W9AKOKIVWxyYW/Mvkkife2SpJPZu5GtXIWnVkDC+ejrO4dMglfKwwwmuZh8+0hIkEFQ1aRn4g5zt
VM/szSAQwWHNMNTzew7pVtuR/7aM+2bArw6PqaUkWLNL/0rNTAc7GtFjd7IOXAppJMiwQO1YboQM
hGxMPmgIRKC+lwYry0v9PB/oHyWgVlpAWnHNETjPyEHmTBawe/YgKjloGp+BAHNg9Ua2e/zeBBEe
3jat4e7N84ui/ghnMp1lcWxsUk9kEgLqO2YJo1NDaAzMjnx/vwB0/GP7AsFeLKjgKfqTj//mUiob
DTDbMc7nX6VLaeJxMbFLRHuvLZlNtv1LXgsWcPgnFvRRp6jqQ8Sj1kckW1KR2mKif6I3KWgzf71q
PXL0S8CUE7SrDKb8L2+LoGVfRn9+cMyoWNHFTK4m/dHBsoRqPDuWBscXR5OLPjI74RNhqpVxsPmY
fdKsqBG4hbMnkoToAK16iZrnPg6m3cc/MMdqfn80QXjmhxYntDxkW7aIGWnWwvlHXKevLzPJj8+h
IcIsUibE4YU/BYTIFsjxRnjhzn1jvsNH8WodYpG9mTczitZkwcsEeQOoAIyqEfqtgYcnuPq1y0Q2
J1It/T3x1A32s9AD10TTTn+w6n4nsBX5i/3oLoErd+IsyIq2E/nVvTOTHLzvYuJkH17/4YSpgIdV
oNcExuz0RedM8R6Y60DfOTddMRJBKJnIC3FFHkE+rWiFPfs25OExbHVEBjJQWrUeNH95luVXzqWy
l7N8vMc6MsyQRc37C039crhCgnMhSZGdfVRAukGjfxYbrEZvOMi/zSybESE2dF1BHb1OqI5PytkD
B/CvGTOWl1Q0+O+PIz4OnvhoN7MCoJAxo+dD+Ee1gD/f3bFZHnMV7ZObY2iAy55LCsH0fmvWjGQX
ZI36B+KpghOUDbRr4FUok00BlKiGlLhXPjeLKrkzbWDncBw2e67GOvohBEnfVOVlPWngjnNfc1Be
GlH8tF6t9VuqgPOuK+IBeI9TiUHynLUjfZ6jhLy7ueR9TTnh3Gx9isabueIKvL8Utd8I/PP7JSak
AjoXQu/HXW/b4GGRLYxuF1m637NX1dDnuM9ayqnOX0pd0mknBGUULZuS9Es0ey5tTxS/wdEfuovU
i6f4LUB1PEFb1dVbpIt7LAKj3k1ebfDXW2VPJxABRtuk3NlGaGSwWJ98WxWctRvIsEaTQpL0p8pH
S3EWKa1NFilnfXj1Qj8/Ln30JYxit0EbL0kPPTPVYD7ifTx5/F58/DYv9kviiHFN9rkfyljLh1nt
pi9F0VhEiJZdcd83XcW4mplISuqn4fsYI7Le9VbH2gEDGEUOqB4eDhG+fTQzFZaz2Bvs+boTmU6I
aJtPisnsC2ocJL5SeOBfVU0CXjjGOkQLlxFe3/2gMkFMuipzr2WgN+1eIyZ6fHm9W0usJdq6yBzE
D/FM8jnDNmkvAUZakVydqZSNRMdbMcPp+y/CD+j7cmzQY8FPQk5NuqxGnzgFrXLySHrJ3HLXyMMy
j3Xp6BthIWDxeZxnBjaf6vYAT6TlFkysss1XdiNXOPN85ZyCPmGs+C+70OtcLFbXrgq8umtx6VL6
WGl6pAbejbqZxUemPTEQjEqbFWkEarZKRnDb9YlXR6zbOUZZHrrg0H6EqNP5Tnz6ASuGeb18dOlM
BInYpV5OZVloLe9S3OcTKbKwZeevCTAXgUH1m+BwG0prAr3O1lSoRbQY5/VYKezpcdsQ8kr9C/sG
pKj5QK5FdtQKMfj4hPgW+WW3uoGFZ5cWABVv+hVgbvrCJHSZgIcHv6l+sBjkL073DbldBYoktc++
phZsxrGtM97wpGXGeKccxQ+oigJLjm+4viC0q4AURjjeueHZCf2NosafcvVPl1rDG298rHh5iCbL
3mon0bskn0fgEe8JDuThn9tLx5y5hCesogXgXLD1UpOfYadqNxoQnZOGN+o7pJu1WUeIEGrAZ72B
oI5WHdo8wU5qnB26L5BzOodw5elPXbdVBj3SxiV2KstJyZyxL63lT4kusQmWNDGT8X1vWNalTWaK
SAZ+5JF7Uri7IDIL57bQ0/VEZxe0AOyHnjPAOECHrDdy9ezsukYJ1KHxGCeexoKg4vTOh0i0xuWy
/LWiSJ8xqxx6LzX5hei45U7q6e2ooFweZXmO2NdOxqpYQwItZPxB9Et667AZROvKLamcp2YDoSc/
+O6HuIO4m62eUq4BV2ILfRKltlKbXPyurPFyur+8RFke+iJbu1jrQwrvhzG8ZJOXTO8oshqYpQPH
7zAnpbYo+xmkhnSMmSCh0KCgw6eXFYEOp3m5IKUsG8aIl139n/6n8aHrBd7h4RUPcBhXLYIzliKu
vI2oYUEyXP7Ac+eiLNU1uj8Ztp9TQdTNBZasALowdHrwZ5GVHIdSnqwMSdN82JwclwwrymWFdiVD
tuR+y8VaLSHtWM27TQz60FfJfC6OUQHMRUeEl6E2hUPlxl43lPyRla0sIly+B97V1IFtObfIqJGs
5qARrw+HIOTY6/BJYAr6OsqGoEWcMAPzLHdBEv65ryYWBybyV6Y7sa7/MelkvfQtWh1jj9tGQeXk
qmDzFHuS8EWVKsP+BjfvKo72UVqAjBk8XCpi3QIekOBrWohSSXliLWYpcUIFm4j0p3BFMwnAcn2P
qUZGdz0Fj7jg3gW2Gvrsi07Dgd4okrtgyclwOXPtm3NF7psU2NoHP81DmU8l4+/ro7f1yeW1WM/u
5Jzp7HGanm3yYe7aVjgfw1XkEzAfuyPOPgsqxSZD79oCEF8ABp3/SYUGNCp9CN5O76FyHLq5vjWw
he+rdoJb/Tol7VSANMbdl4t4ggpibWZD3eTVt2ki8T7N4wQqnQj6uTVn6xTtPmz/Vn0fsqLoo+4o
4JkXKeG8k1NvAVsK1Wbmpi8tDgQqX82Cj5b0hVuWVzjgTQ0esCVdH19T5nOicvlcRDdwoAPzpBlt
ysJMC83XUOcxc+WMd3iCaAIn8VkUZyrd204zCvUYR9ARAzrhNoFiX8EgbY5cZt5Y4uzSpuDPhAqF
Ew7eAAKI6yroGn88qaHbKeA51H5cHydDTqd6eR5N1e4sz9Ydlf9ny+tN3wgW4QN620LkLS84RRTm
wgiNBzIk18Mox9zDi7mkTd6IgyynWYo+EoRU2NOfLHqFw6FkY3yf7IZym42gD3OLQ4WvCl4Tv0kK
AIuUtgAIT22bmmBSaOuSEdHu7oE3CNucAjTm5HogaGp9Ih1cX8lzHhsTUaHiOvSCAPU/IaRXt9Sf
aMQGTIPKi6MiDn9J1wu7Ftuwylffc/JNvi/FDJPc34gNTEjVcT3POXqrhY+KH1rrNJf4Uxof3Fj9
xhxjp9tyml6NXeTmGeUqIcdvR4dKWsL1P/jRJp03A0zEqpBiODjc53eSh7HnkByD+EO4Hesh9EdG
1fUxN0bVh31Ln3IGjdoa6eJ0HNc3MX65pEtQ66d7dQROroaJcg82/pKwlZI5PVMw6nDMy/p8AT4k
HUlg8ecuoiL0DxKxDWCXR9yxwz0uWpezmO7VkTjxvY1SNL5u3jY3Pzg+WOoVl5Pp5LnquWnxfFp2
qLdoedu+DZfSsC8Cu0xa/ncfI+521UjAdr8udOl5brl8r9Nfv08Oi4YDeffHs5kseknWP+HeQz/1
d3U1Dn7lpt21wcvEuRIKMgw3I3sVMUy0fjHbOnGtgVDRdyaxXbpRLSC6XdefQJPmGLzcET2NdapS
qH5ByBEfRnXwc2wxVw41piYuRUCvDTE28hR7wBumg4spvpYT39hr8Ljyr2hIFrHvY/oA1DqEIQ7U
NDZpuXimIzzl/ejNVr7V8yfLw0fH51245PByngvr07nqiIG4yad9E5FbxU1M2yk3FpNsHeGtN4gz
wCz5OUXSJRMqNtYGkBZH8oqU3rTzQUk35MRdrtEZiw0JmVnOWQ+5pJh99astdsuvaeAqm/rGV+CD
hFxsXjzcGDRUtwzZk3DQcu8GbXn+h64HwWQrQQptHnfuI9uT+qq1QPmKgKmF4LRQT0CQH46eQqL2
XAfdGYOZffTVcpRjCATgzNF9OR+d6hVI2FXPsD/ivqWzodA2HnzzcHRc6ijjesI8JKa+NmRXsVwm
DpbeZA5ZtzJVGo9jsH7ZqaJWQkYWfokRjqjwEOgQD1mwmIyCFrAk1/E3ly8G+cljSbn9u9baYFiK
th5nSWrProB0ET+AnM/1rZ7sclaaK3A/0g2mZ2J1zRrWEnM9mJOBbRNRFyy4+yTrY9oppihyRMIi
5Pvu06MxHFmuBXn8R+s5Y9pW+E7C/CYeT57nX2tv16RWN2X8r6xKohlbvimGr1svmOXiXJenHhSH
Dmd2x8RQJ9OVLw42gZOoAE33mz/Js8oDjyuZoGwPoBpf9X5cDxwcxGtamJqBKktVaFPwlJvmDQyu
tQXYew6qmIzQ4HnQ6VrhvxXZ1sZ6bePETKbaQh/5ZdoFI0VqCwyvU7ScicOJrGzSRd0ld0AJe0ui
Uf6OuezFUXeEIJiL499EyEUZud3J1b1E/PDALRk2Vr1KaX9j2WoiC9d7ZwBNZzzrMxSArQaegueM
RjsumpcOn0fXqX3uShH4UyILd9xR91GXwi/my0EhyrNhw0lvtuvC4CtRWbxR+LtoWB/aV0A5nG1O
vQ6EZTUfJ/nV9ursq7RpzPDEPWPKTqi4gfE5r/xs19yL/uCQd5mIYVXW6xxU+iUALXp/6Bkzvsvj
Ta1y/O7zyjXCSgPZ25DPYmsTIkglXHzXaPi5cLIz/4uKf7wW+nwaKxrIdKjg+L7ZltjvmbjJmYmQ
tW5F7rnrcEGhqY/e9TdaDLzsj+ORzB/WZ7spw5v7QslMp9WFerwnK3Z2Vh3zKTvY7i6AqYKEHrjY
y9SmkDDiy8+lHw5ZlknDkIDwSGAIzgOwATiSjwxf4AtJL0OcWogqf1qSGJYNzT8tJ+ZJechirzYK
Xb9OmzxNda0EqWjozWcgOWJEOZ6dEtK0XbNG4e/kO2/cM67uzQq6L/DyQzQXfAXpoe6Ve99tR/ET
skBUO7Sx73yGqA1iI+AVqjvCAEBtJ09yV8EOJ3npdTCdkZS/9skmalX1+u2Y/HziAvY504AKqLHl
RyQxztImlcUAEbihs8zQrW+T3WrZOJCwiuBrfpWmwvu88vzFlFr60g5dqfANL9gxyn+z50IMpyvY
AAsX84lGMSwiVqWPBOAdV8sFlxzX7ZRzpYu31mQpTW1IunSH6fmMUDoFrmwb+S7Bwpa50wcztxwI
vPoDf/usBY0kOJv88rsaizN6oge9CVHWdJ86isoCoxrtkaGTA3MquPR2ZP9fl2MwcqrIkigVed3o
Rhcp2dN4IhFh4COodOCuZEvstVEZM2PQpDZ/QkDNjwOecV6hjuwJO/DbPMkE+Cv3RPLE1Mj/gFHX
+bEPGFbYJ9iPr3DSUnmeuMIexw+lGSYQ7niFXsTlNVuhPkAWc0gxQ5T/LYOZ1+czioy1JoUy2k0E
QPXMIjGt1g51aBPbMizKScdifRff5xopBDwNcz6cm9CnGcfTeODNFbC2DwF2+qaTSChTMn3dPs8/
f4sSLMVu8/Lo778cPxGfU7oBMZSoJIypWzjPwaqH27jhq9sjEjqEwutN7qJldAPoQbtT2dmFum05
KViU7g+NWE/EriAQDywZrV91c3FznpamGfZdVo4FKgAlqjo1+ARNbJbARSQRq3SO5JMVswC1zxMh
CjrMpYO2szDw1r/3zRY+fmPhs2EY4aCl1+nSZ2tn0dQGH8vUC0qSAycPcnPlRdL7U4pitldBkAxc
6njoTlI1NmPyTlf36mF+UnXrt/0vXweawm1ZG1ozmi4AsOGrrOC0ffc6K4jOQvRysTQDCygpnqc6
noJvbLiI8c2PbygvQE8nLFSQE49YIujuxihYaV9Zm0+Oy7mGck6aKlIhOWtDUqoRBX/zCb7zgXOV
SQMMipI4+u3GHAF1XGrKHSabQqqY0ZhlU0bpsi/IxAYlbBfXylRe1Q4y8OEQsnRpKE9U2atJWrc9
PdeiMyGL7TDh9MYOKjrhX23HOxJ+1USedQwjnoGHzhqOhWNqBWhw/bEShCSn9Qn065RrsXeD4EGl
xOlDqQNFKrSrviZEwLMFAt0jVcWz/bwlfj3T0BTWv30O/a+cVTSQ7bNThKhTWpqH7hFG/MQ8sajd
0EgzsBzQULNMa5hWfGizZYWe5LZ2MjDte/qT/so0fjqEdAyQd81PovEsLeeImfVCRKulb7ZOZGw/
B69hn9q+Azo9FlQjRfVvlDdv4K1LqBy5ptfxOdxTzhKfOqF31hFWipmdWPamQeZeeTfDfF/vJZeg
smxCmktWrXzlVvCVmND0Wa7jpTKXMaZGICH1GX7ORvqN4bJafoSy1r839riOrB73fOqPwP1CsCf8
ataejAfKv32BwuMvPKJiPccX6C9WQIT8XIMykx4lurBU0Kfp8t1xd2CREfPSwCqCpfEJRPDxsL1h
51qZ3h46ce4pOrPg+CuNucd51gMwcxxJscnyPCYytKT8oLbKqyJlf3zDJnjrlq39D1tXvS7IyNLn
yQQ13rMXjp/gW2HtBEwVVXJ8D2TZmck4D7XidM2PsGLWHjCPUKamZG52e9VV7dA2BFtfzc+fNEqt
2XQ6n00bRdPyFiZ237zE5fbVr+Tu7StxZMOP/abd3G4163zY0kBU7pN9rfbs6qKJjUxQFDz7rhiw
WBWev9teqwHWo+n6lYU1LTlrauVQ90zh7VXofSAtWGvjBgrh/jdj0yXxVh+AkWwi5w1BOW5xKKwf
7SX4f0a2RzwtLgyUUHZtKqc2NjwBxxrKLC/WmER/u1E45OEPB1XFRrO/I2XtaiLQzFdrK/wvztJR
qs7XObGyqsUXyC34Fj9nl0avsFE+yLv0J/+Vj8DJ/rzvSn9KPK2IEre9ISeaGYlYcYaSlADro7kS
xwLOGcSGEa9bnP6exsWzfwA/4Nrv0tW+cfkRxmOohqlEjuzgi1BXkm8urQK46Mk0D5QRSUeG1KPO
T427qYw/tjG8yOmRtpntDJW3lmjt6IVFoxGTMdCpIiEdBWBYOmw73urtT2cPy9YNicESZ9t9KhgV
1ZL0n5Da7sh+2vtocV3iu3M82aQ9a3X8VcLEaRRyiIozAJz5dXwAGy3s23DU/CvQYWhMB9P07FE8
yAuR5cgMOpXcfCRj6gp3AEFdXX6q1x5MitijLfxuQyoQziltgbmmJ9gRrcnFRlK4RG4qnR0MtTS2
bbb7xwOA0EXJJEAYtBOqGel9THCIjVyRfhHfSEVDn7tM0ESagEAKUNQ9v5+Xgj+gaB+sqdRdGqnP
lX+TD0msZ0jxLQc/4g6jV95cuLoRvRzxZQPkZHi8EMxTqgWOlKUOOJP3pkdIb1Mhvj/fr27joJ7y
Dy+nz+oiYc9IvMnwJbM5JqieGUVySQ64soyKNzvHxtLVH8w0/sHJp2L6NGo0hiKMZkTB8P+zKu98
fnXhQVXjtVAuPvaWYWdTFsQJeg96zKxzkLfeoqAU+BD+nICj1MjpWB6K+w/gOI/Yy+nNhJ64i2Fr
Hr9mUvxS5cOyAZMA0ze79NFSklj3h6VkFi7qdgG+GiIG7aY7xhsTwsmLWrBsCg1Aa/Yhc9qNQpKB
BLRvLwNqbUuCRCrzAZCvTl02YPxdp/YnfUeASGCdtpjUnB/MrPoY2LDZmVt5iDh69eVxPQ4GDuN1
i8iuWDLaae2QqBmyoKNvfejend3VzctcpZ4tfLFmliqrKDEgLzQ0PrFu56OCaXHUevcWrSFA3cnP
MV0M3GoiP9StfLJ+nSgZi4HC9ds0OYHBKAXMGjk1gmXHSkfymI2Bygui3356Pb0+CIzxPeFgF3E9
Cwsy0cfNomZ659BeNeWRTmR+C4r8fJA2ZC+lFpnXgxztIUH7C2buABfZ4oecrepDAa6fXrFCkp9D
dXDgfKa/jBBLgqiBTol5W3pwA9yEHfHqgMiJ7hkY9Mlt5dRn9z6G3pmYrUozZS+dHcVVqG6wAnAb
7Qun5KluVfFcDR1n0sgK0YUq/sgj49cbUINdiZYk8JnPbNP1a/OT0KRyb+6EWXyJIfnongPLCVRC
DiOlRtQlPNLUb5/BkVlY3Uo3RHSBKRIIFKXvKX6UM6hUPugFgOmVXO/qalVyZhAoNM3gEAIPagN2
VFDCertPTXedFhrsR7/ewQ3WBoKowgTuYEQUSZgnJH1UUolhadT2bjhk0fN8kW55Jz67+UDR/LWx
GZbawTKzH+qc+V+8YTnNgNKuWAlcqMiMCKB2jIfZMP4WP0T1l9Ltzzq/zFQUQB90/ZZIqnOhOppW
vEwB3B5bcVKf7VkEYCD9GkdGcsuzN3USBqXONI6xle5K/PTWg8zY1Ww/asCAr4xMXtVAKrKrnUP9
VHKtr8VPzeKyWB7Vf8Zk2+kCLhjozwJHR7sxYbWQxkGmKgZFAD3A/q57XGZ292M2lzJg480mDEEj
ioht4+aDea1E04/3rajrERwoPNYy7nC4JWZo9nvcFLZf9hBJPOmmBEmeJRqAqZx21U3PgxxlmVYq
LLtPXgt8aN0pKpto7zqX4Kf0K/mgJHkAK0J+blYNSxcsXrSTcqzHhrSotczQbRNTLHpc6ufS75Wv
XR+xKNcXMUGX2G8G24+t1fNCgmpBeyjC15mWgSotovOajuSiDwiXk2A0DeGOLSrk15ZgYoe/ZONf
jqe/fSRCw8w9ee96eEZvnE4tq0lwH1gdZ1zv0DCrxPFk0di9K/H9hDrP0dq2hTstz+qjTe2ZGYSf
QTwla2W8fj2OA1LJG0ySrwkJWBrZmgQcXp7ykTwLWcGoB9MX9ar+MWSjJrYrs/tZ82e8AoXgDM14
0xfD8HkUKX8YCqkV/+hkxU4rd3UEZWmkV06DdYTid/eaJZosjLh9flcwXOhB48uLmTclt8a273rW
TEDl4ab+TwhTGAWYVw8f05Egqr2t58qOt740YSOJHwwtPhSK/rLgq9hjZu+33sbj3RQ9rBhooF6I
1jFVktYSs9YGkHp3OzBh+Dwh1E8watbKG8SDfysKmxOQUcwgV3QU6PHdHqwlpD3bqyne3SOxTKbQ
HCk7GhN6qEOscgI2vKS1hBsfLw0yW5B9a1SMZ1hKs4b69l6rc1eeO45TJftRPrdAFgjA4VtvNmA+
rY7PlvGrAsXNgbguen4mCsfGfcrzRYEczLRukWXeygsy+IlKdMFb/+fjyparql93trUQ9e289REd
FI/aLjWHvRPbRHGZOEbkfW0uDJpnipc01Y1G/pPJeg661D25KSeTe+Z7Xmq9z31+1vdk1fvwHPG6
WeWNX8TJhsKp/sx1Y71Ogy1AiRsN/Eweq9JwaICSYUj3uOdiw+DpGcm7T/PaWINB9qktMPb8x5+1
dikBRTwT4qClnL/00GE42Cpiok0zQonVRTJFNEdTNVNospxG5ulLvPnB2RTbIzOsclSbFfffcjvb
gB+tOHeByaoAMzFOMJPhNkOgHsfVQrDgsvXgIx5FFdyL9NYxPtYrEvyq88EIWovIQA4N+xmwk4Z+
GrXovNKQiAS3eiD68P+Co2NDMXkYKEj6IOPo+BVJIXyS+hjt3ptzfRSw8/G0mVBlfV7EKZmxmeL8
WQIFeRs20I7nQfWpVK+viIKVjYSZtgaK2HGd+3TH+b81CG3BvkCNfFI6PKEfXSSjKKLW/yK9YShR
ffLMF86ApuMYjZaw2DTaxIlRWE2vYtnZBwT6CVhrwcZGI+4HyafaKUeZleJMmC8jarVmrT3AV4uS
fa2Abd59Kg7oOSMZo6lcwXlS00xZPzqI+UEvtXT73CtQuFStQkA3nlB8hJhB1PV1fKiUHK3p5Nqt
R5gCUvoFofVPHmNc0BkVtNJ6yGBsM/zKPk6lVxr4vj30ONwxHQ2lhUHWrSnhgtrSgjxGTpB8YOlJ
L2toPRUeIQA9oXdxWu9ySgiphJ91iXGlYNRjK6lDmf0h26zkLNnRptLnOi76gHBPqMrMAVtFwJ0m
IlQNpNtRaTFJ9Y6tzQsx4wbS1ssV1qZOnDDI0nm0lfOssqH3Gv/kIv5o+6ExVfMpZ5+HYUMGZvHq
llciOathuiY3BfkqOsFhiIqz2+/b6iBbK848K21abm7R+ZizJbffEOG8eNtdE4V/hKCyjTmFDokC
qbmRQ5erU1PCCkhQosbpqaBNb82grqkkPT+MguWdGMqHybzWZGBSD8k3QauOCdWdu96rbfwm2+73
PbWnTaUFpA4bg+n5Sl1yJIp6HpF+hutWKH53rzmwZz+odDMHl+e7g2ZWF+7bkOBNy0QsrOnQo8YM
v3qb08IRVvqpIbdIXPcrs0Py/Pzt1whacK82/wcDdRC6KEbc7QtgTtva7egjQQJQY5Yh9DB4CMCZ
vkwtDQdPglFLjDsI66TqbnzuPWGH0/70oUs1QW+ShBqYOHI1egFT0HIN2OBwufXYGCDEe+0F2tZ4
mH7Ekrwzl6t1QQSUkwuVliy5+9LUVjdZEnLx4UQP5f4R12d83nk2rxJ1d6ZSVSIBYdcYCngcmuzf
sL2mpt75ECe1XTkKJhc+1qGrZrAkkQ0WyTbGgq4Wsj/kR9x3tEPKTn+fdGNKT0HzEoVmGmkYKxbm
dKLLJE1hRU7QphqAw9gnaBmpOTBOSyK2kRaEWmJjcToODY7P6bQ3BbtH0EFUluwwTcLwWBrHhCCC
ZbAV3T0mPuP6roP9u97BpmFmksxQNna37Hr4ZnH3KtQjDHhnsSF5Yog4NuY0rTP0rwYScBeSIorD
aZSvTYMibI2ccINdQyH6DVNoVqIW1vtdEWWvMybf3Vq+D04nRSGlZjHUL+zfQFJmCYSdq3Ltmyw0
Ppx9xjkSVpkqnVe/LiSlqkJbl+jzaGI+yliIQOyAhgHr+JLtrFyxovQuddVlNIRw2+IW0T13ouNy
CzquZDhk7gTRI/91H7x05pKY/VKWA5C3BSWy855sBTYSdDfX9q75sbQyCo+d28xeRHtniDpCVm+/
St+32D8YidKOH1nCE+IcSB3YMrV8qPflngHOfKb+JJk4Uogu+N43dYzwf0QfwGkFGZiZwqV9vOyW
wkQdtZcD+7nGWswqvohwIudFomZVcvTnIdYocC2jXxHRIuI4BRhPWt+dZ1B7ZKLiex2kshT+oTIO
bZTGYqF3s5L6jPra0sBDWEci8LNtKo9EzG6KAvJcT2J+2kswuOZrTWlaF/SfzbASaYlgWILJKCX3
DXqWJpyWjyB/v8vyo9Y+H0gmTQR81KV5EQne4f5e1xZqjZo0Bvgim05k6GRwGbssEOjUr9mxbjIs
hSy9WvvBSywQ8Shq9IhLRYIV12Avvo8IWrSEbj8dzK5kXTB3x7+VabmVHsiQoN83Zysqhz10OeGm
AMfyxC1H2t87g5sL9iB+vfxLU77d7KBR3bFDVn8OhFddVPKJA7wvoVTP18Dbd/WagluurGlry4E3
Hty+LgidU0oQzHdSxsIHt/trVEVt95zeJePzqrAnjMat3E+sjl6ARx/VPcKq9Uu9HzP7fpx54VYc
btXmTlgUAbhsOvz9tadayGdoY1U3RKsxtEDiw/a9nuYzti2NfXbFp8Q2Twvr9TM6KtiPM4He+kid
xje5gpowCWhWiLlEek9IP2k/0ewXj+Aj5fT/NMWNhP7HiP3JTR5515rvpOMW+UMrqk47LbjbVA9v
hbUqop305hf8sKV72h1N9ZC+nmicORqz3KVeif32SMIRSRV5jUxPBQioauWT9uoEl5Iyq9FW61ly
rXqE3QscHsWJOTgvCQ43qGpkXEPb2La4TFpoNMIy+IvQKAhgxRmLTMK0Y+UMUuCB7TkxqilDuXb5
LxdJvFOXFLLI5pCkzRZZqx+3mrGFBUsXDnkroHy/BfEYwhDQUJu7lsu1LqbbuFr7+3CEWO3SgMtf
r6GKqmudiSMFH0O1Es3kZMuu3KoZtWSvkOJ8h4gRfQDFy/VEyDQqwpSNNr4LSkyDKyxYgPFU36s3
+eIF45PP0dYCVc5HeH8xyScOvxQz/S33/KaGYygIC5dcoxOfoKfs3fv8VAXUndywARqu6L6mlF8k
p5aT0YEOstIaIbDFL5IgWVtFrJLVLaKd8gLNLk7FIG57IafBSHzLMwiPW0p4Zthik7nK2EGtwQPw
VPLaEM/3Fw2kbfuQkFvOL4n6+1D/YKpg53ymbzV8gmZbcqcmpn87kxjmbjKXnw1xu81u5Cfcs7g0
uCCQg2CbnqVnQyZ+SdnrYIeXkrnboTkzPQtFAbYDlVG6JflNTXvvK+y7MGqZOdn/e3CPCTkXb45t
lyodEbau737gH9dT5bnxtQpX4nF7dHfRmqa3TWVISahc4x1v+MxkrfP2TVqxjyLWah3JmcwWxrkf
3sad+6a4Tuw3gLtodFA0rD+XTaCG1LFc5zMECm1GfplbkqAITccKP9ZdDtcTiRuKuxhbs7Dx3NNv
rTLD0LE61wQKTDF0c5UpnmcLRjHD8IJ74uL3eAzVt1FRqd6jiAMrR5gy0kJIRQEQtgTMXM+4/509
8IpyLm/+sH3hG7kgmOdQhqV69a8QPdvcwGYuyZMfb9BS+RAUR8Jksb4AuM0v+EKvNyfWj2eFW9SB
obisfE7t7SX7QqEV621mRAYVBCC2NqvFaSAHgJi+7NnfKZtbK7j1DZ436jgDanS8jBtJY5vWCAGL
3+KpdfEnLTQ7ShEfmdjfyAq/WtYKbdAeM1bwV6qVj82Rj6GXcNB9SQelBNvzYkyh/C3vbyNaUtLo
e4RfPhFETGzG2X0BVGsR37FkarELCk0SdhY5OSNCz5qgk5Tln/ba+sn2Mm09zxUYyr5YsJclPouW
rYc1QNFoRLS469Ms/lagncfervfR4s1uTFU2DPAa/JM29jEhfJa3+vflSx8YZFlB1dXjgmbTwEoh
yfhHwWMZAVUWNBnXKHfgLVhDBr8vnV7DBq3Fnd8tLNR9X3UwWzmW46Nt2gpc7nEFavNqqHvFPmia
E2D9SKRLe2ZRaQqdf1CF/lstTLtLEEOWKBnrj8vmbLkpBnc96TKMQOMmrj99fPT1DvgDLWOabBZ8
azom0GpH8iUUxd10yj5vrz5b3YTxy1H3frM+kDBi/iNzu9WaEeRdJkz863iA0IGZqrW48AAF2ZGk
8QhhCd8Nbz8YlqxC2GE8m2u8AjL5D+DozUScCWWWedDRnxAW8lqecAL0IQ/0tWJfRagmjlOUSmj4
io5KEEwRs6ixAAXkdCA0oCAhNgrgCW4Ppm0w8vTbRzwyVv0qxyceMxo4vlkeeZgNEeIHu+OBPRcc
YW57iCQ59jEY334/tD64ZJTTIkuTsWVHVBduZS4wcoJBYjarbN/a3BgrVd2PD2MTBAvKSi7+MgZs
2odWvK1+BKP8HH3CYhgafg22dWamxfDKMHkaepOSFkN/APjUApbJBP1J2bvfKiJ2av3i6IHKFFFv
XVVKzFisoPC3oUafwwKnbsuYq9rYuwYhchQvI9o+u47Pxno9KQjFp/2Vdfbx65woA9ldm34BRo+z
K3jgWVntkiq5/CLsRXFS5+qyde1MLQ56bupKv3W8psDFsKHlZZgH6meNKU7tjaIchtmdD/69SRjF
hcttx5AIpJdCLLwPG6mZi3H2y/9mu67rRAIqk7OInnJCjAR78vnU3hAFc6mZQzF+szgtbyewZ/ES
sdUFvuPidyxFVZG7/P+MV9ooGDuRSNC/RZFtcVniJM5tH2yqn4ja2JyEPxC8f+uV2tZ2EryJjm+3
IwDfgc0GULXJbI2lCCJ2JaWVr2/CyxUcQKIOYOmJplFf8GXWvoJAJGNF9KFvAlIoqARRy49XpMsc
gUswsrz6ykZGb+k/7griuwsIxg9b8Sdl5kVDSZdNWdDQZEqN7dtkBpZHfG1PxF5hWuBba/RhbAa5
GJUcDzm8+eax/83Su7QYZK3mbQVLypZDec3JuQVsL59veF92UvD84pgr8VSPKO/Qf6zwWvLx55ml
g0qcN4C8RyPBj9gUztsj+LtfadRQxX2p4ddeSHdKZwMpslwS8o2poJv2iuaQAAgo9W7jwIHKylPR
A6esoDiZDq2ywQcGGxq7QMFx4Sapib/TwLXwDw7NbHBixyGyuePDqfCkxEFuoQYnVbycCpjwIgnp
UDVnLauHLNgeWF1ANRgZuC7MbMlyxr+oH/JReZrjkZGsQZi9ftXnaDNJLYGr83Px/UryD8WS+XxC
DdgfAw0QlqsDgtlMkHwDX74S7zxypOlv9c/nJxkAIKCO7SgFdPR0jUVPuoUifmGtsltrq/8xJ2Kb
EC6BFITKKuTEFiIyjeq7LzdXAr+ePVWfMvzNP3qP8YXHPX9M7H/Bs5Fnwso+xE9ms2JPrEoqLxXT
ds6jD2hLvDPDgHSdCD7UULUOAmyyxL9CejCz8fWqTIqB3T98vA9Q3oFM3ObWR/ChWbnHBFbKtaW9
u0z5L+BTVZe+hLXph9ZnC1pS6SJZZfwtStsG5Mr+Aj3SwwR5C9TsC2H54w2Gq//iXeior5wLQysD
s3vEfrLDawHIvOHbfWwZbbl8vGvaZ1b2gG9G/Ylhpng6qUNLmlN6tReJv9Uf8NoCHSjlvvRp0MAk
zzJkV4+MXCe6DWJhEWWMmZz/zSruUGAkF1sk5yhiLTqZRMq2S+zPxsD0VXIHiPTPwAQ4IPLwJpoi
17UwZrMlngq730oE3i6/iLLCHzeLLuVBlyOJsXqZdbUm6a4qzKtgxvyS0ZNhWZKKayCxKfcgLSmw
uSDTz1d2iGqXNDyAh3oGDxKYbRI8LB6vrND3bQ74NH9ru6kVeBQ/Om0/O3rd//z2Ee5hbLGfHoAE
kiY3ZISoLh0AKCXWsEqy8+3oUQZ0nUdh4bP5nH+EM4mbsPH/FeICliZKkLT2OvgAzgObNaVqqXf2
cVH8R71FeG4d1k+XgUhoegmG/7glwvN9pe6hSVDe0s1Ybfj3mfzwzn21eRtiiADO4B1b3E6gydmc
4JIK9s5KwoNItXT8hbJ0CHutsPN6TQr536PIbBFGUxQ3Ve5XzDB09rpjtPQSjO8I14vXj5hTHlnk
8j4arjYAAPm18R/0VCGrOiVKOuswRggr+ZBQ1yk1ev1Azej8Tf2/ISh9H84A3RSMn9l813eatgIy
iV++jAbWybfDiEDl81z04nUt2R1gBxolmiwbCfqz9dC0rDVq0QPil5wy+b0HWryOqNpxrzeEBYWK
eoDaLIKNqYi0hgU5v8kWExFSdGinIcJktpS/d+RuyaVFuE3PbV7LwshhBGnf7UvqsWJlpaNEiJp7
3k9FZj4M2hU5cfPvyZ+Yghwe+ncOCgOOfv126vhcUO8dj9YKZaEHc0+rPdtSJ8jdpzu+SCt+09Yb
sO2eb6fL8NOj3zzfyO8tpLHVpqSUP2M4+sEQqRrG1hkBr/2JBZbCRrj2PL8YuWp14h161k1oMHDh
SiZUbdu7fqcZu92GjxbnqhkLtslfPiVtywiX/LaFFyYqF3ye6zMKiZw20ebibSMIQw0W0wbrYqN3
CvQOeJ7TMDqzEh7qs6kO3R8+i9eTax1LxDyD//tp3DDVUpHdIDlA4Dvy4l+RYi5Sf97yr98dW1xo
QDQjOUuIyq8v8/uqX7DxdRlTiGraMMJkqDC48QoaRYDuAu6IaQoLJjHxvmkfc4p5/VcRQS3yJCN6
9f7teilBnePhWDUsXTuKaakySRiqdAhYrkabbMpnpC0o4kAv13Lu18NUf3yZZ6bB2ijjWkcLYyKg
WLkCrc790zXmfzllP973UzgCho41Vwz2Nk+dkUGRxmDa6u1S30BNGNidF/CcE+sMPN86pXceC8xf
Fd9YwE0SJPbt5Jlh8ZfezJx+qtLDyyaPwOD5Ie7rIg7Cdy+huhNielPnUKq0deB4beMBqhpVAl2v
CK6DToeEpSQCgiduK6M+QNbk2Bl6s8NrM2f6oA/A5fsDSEZWAILL/krAJOVCDbhTm6pjARks4+Lh
WUpDoGdBfHo4iNZICn6IPBkE1iSBBRDkJT8rq8g1RQykdK8yM5+08oRUi5E0uS7PVAG27/Kwc7lK
PL38D/+sEdFwoopfl7iLQHSVmMdlbCloD+B+o+TnzWba8bzrWMEPB7v9ZSOhyxhaJ9q1TLxitQvF
oKSX1IZyduLTgqEE2sBQxJfnvoviMqC3S8KDjMLyjRIGd5+c5kxQLpJ75GxKEHLAhzUNQ4RQfKJH
L+1Exicc1s7tblutYt/17Gl9AU+L71KRPRSiNo1RiL3+7yRszcvQKOz+Kmqwn1ONTclb5Q9sy0dW
gqvWSEHRpdlenzGm2gGkUOUcrphj/wgiDbLLD9NRN2uN4Rsk2MxQGZf5AH/7zO6xocvyuktuSDJ6
1PfWBRV5WAZghhargN01fcno9ogUxVklOSSGhJMecWT6MF3tefNJ+kEj9vYGQ27PDpv16nukgdle
g5BG9iv3MLr+O5PEVr43w4RxQ9a3RJ79bDH8v4xckcaFgKi6rMemWNsnezZPVUWf74VHz4avWu4i
oy+qSIUsdoQGiSypsb64vdRtekp0NhZWWhKtQPO02NR3XcTtWDxeupWf1lsqWyv91LkiZ5Pz0zx0
oaVGnHfgLD6sTsukTnI80fdQbAEcJAXS8TDTd9olWJ99ZHM0OlgtJrS+To4NX0v2gFEnPbEsZ349
N2m5KhmIb+fSWt8eJR3qEFkEqJySQpwABavx7arqkA83bLlhEa9m0iidnPXtN3g3+9foluuMrKJG
Y1/Rfce9aH05ol9LaEUflg4movd2L9ylo2NNad7XrQP0qXZIFYKRXMQ0zreU6KnikQKKAQKGzRjy
Hql9xU8Its7aWCqfg6PBa3CDONuZZ0BAiTm/UxHxohBszVVNRVTTdeZviD+yQnH9bqh+7h73+77/
resB8iJqpnfUyPykdp9ITlfp/08NnQpF0aHBe/t3dze6IBac8S9it3SBFUVxjXkZzhzquE1ls8UX
sDBCxmmmaCRhpVcbt1m4KyFIRPM8NZZPHuQB7tXteAQxS6Ui/sZgeeFdYm3EcTVrfDBBrkyer4JQ
ONf+AwdOWuxVO41SeMEnqPzANyCtueO33Atu9s3W/tMJIvUxuvEzNsUJNTvly5omSLdnfw7tqKqt
Z4k2tVdDZtaeiuqQs0XRx6ebseY+PrMGdT2HIMeCQOF8tZDt7MNtA46WtVwL1DXLnxZ2sRluuW+A
8kCFQ7HGZphNsIaLBuq8skKC9LcrdkiuTglTPI9orWolgQjF0Q4ZxveLphoATW4YznuD4QNNhtYZ
oFkv0qZM6E5jZqKgjQHxH207NiYQPZE/gC5QK7RknJ2XL5e+3aigxa0TIlk4vNlxRZzsZsLqa0Bz
4nNBL4VdndpOfueteaRa6N30T71FiYokb3g8Ro0fTWg5ANhKwFKW6Zow+25o5399TYdhTPtNW1ZR
WPUWZGzirBdzFp0NNrV3YO2aXeQXvKpP43kfTOR//2yM47FLt43oTfh4Gx0L+gi5y4IsD8Idmdzz
nTaWYxHik9gaUAq7xYg8mzmJrluqP3B20uPVRqo3Q3EN9DDph1Ighe/YVuo6V2jqvkPHXfTQlEcy
WwLLQRdDIXjYWBN91eC+0Ov/d2pRhwdlXkgaGdeckH67y+5rJMVWr+j+NdDO3NMrEvFcTAikvLt1
CxFiVaFxplhBUverqhZhbJeGRYAwkrhtNX7b3sspvBhhgJ+HtLK2qyMomFhIGnNS3MiqDU4bnnQD
vu4olF9HSSj6B9wUe8Ab/sErGCIrT6ERtP9KUhjXA287juFnobsCaf5nYQZyFgNRRyEV1F2X0Obm
o8gswk7BQvl1Yq3gu4xzVmM8SOQ4LKMg2ga3DNuvFODbutabIrw0A3O4z1YtRFomO6i+rxVARgu1
vPWUdgnpURqdxHPL97B5gIVnSidkFAQ5gJguGLQ4m/jKKE4CZyF9z2/pPdcMkwzhABGzv2fdnsVr
PVVMinVnhSvH4cYu/a988uIL8spfCkBU5gj/SEPZ0sK6KtXb+jiCl/ND5tFKSBZfC2mi9POT5acI
wWjx4/E+4khYppPigbHfUUMNe8GIx9XwvEZa8iyPuDzweFolaV0Leb22FVUKmwNGPFxGLmDAEfBZ
ZIjsPIGdgrffaenQaAnH/nTpHLz4QuoY4qsd9GSm9ro3rzLP26MEeldJLugNxkwjv3K5UTLT289c
XdMSqdvoxkoHooEo+W1JZBNGCA5z/PRKblmX6evxgbGy6Q/+UL2iR/+nbduv2Ll6jvDm3s7cyDaI
s2amsDygag1R1wiLaSYiWxbkt+2ScLRkL/5pk05gXGAB5Vlwob6h401hdQMSVTaKN7e9xkgDPXy9
hVz6WYkYtSxdcCBmV3OEyiym8RIaa0/PDukJ5IOuDHT9p//+w/5lRZlohTv3gEAYdpQxJippKqXA
XgHbPmMPA4qnPF9MY+oL66CeWJd2D0LoE46Hx7Sah5ClpTIh2+FaMBAReTVVSDSMOuvCH9aYKCpC
Tzv97zWRs6/DYQQjOa0JndnrvukHjhkTpv4Hq/ELo1cggI/AL4ckpBqqY1IOG0NWof8nb9YAYRTn
9IbQ15wdejuN3+8VHlguwq5wq2BMQV3hyOoeTg6Pzzx050pVv9biYpuHRRCWUEV2OFdIi6FsyPxD
PM1lvUxvDo229QkLgRYwCMLrxKG6t8WSiYkY6cK6GgpFYFSdjyWyw2kb7CHlPJgK4w00DELKwLCB
Yf5mQMBEWeRgd4ZJ3vhWwonjAuLFcX48rxIufRiOqEUfR522v1xbmanfTWGdlv3uQeFbT4sONluX
P3VRXIkUXlIziousxHuRyk9Y47Ow6Rq/kt3CbjhnWW2KxnJmLL5xW098CETM0tm7FJRYREuymqBN
43/5RIDQ9ziwMhBzQJKbsw9zX7c12M/d4mqMKQG9blgBuK1Tbg6GHR7ruZBPefwystfurOI+rwQb
FkTOpnBnYNvMFML5O02uXDZWmZb07W57WFp+hgSFzpdAUZh06gvPJRHbw1efUTM9JoPpSsbNYmVA
pQ8Zd9SqdBDVihwT4M85hnWd2fUSUWl13Y+KYu/4gcXKeD3uX9HoR3KSxKkHlcqIOSyglqGNjPbO
5ZJ+83KnSqQbacdk454U+/GnYyDIxwSShsAuYipPQIKjsJiA7GpL0YqFqUXh/smJzJbqlhsSSP4u
YopaQva7YR1cZDg674Iba/UH3pIsKN4p4BjlFz0f1Q2ybLOcYP72DrRMSTlM2GJS1AZbiziQO9K9
inegs/yEkSGRwoTjXzZbMTTqPDUQ9fcjcDvM36RJ8jh1Tgfm8d37eE6mdjRG3hEIqN3OmoCCbnsY
+rBpS2dR91IV6p5yyhAT89v0BIwW+urZA2qiiopKAjFtKuKthy13jV5iQSW7JZm38VGxuS6KG+QT
MbxdUZ5BGmvfyo7dhJLH3RkiotmzJrm59eHWsAkW3y7O41KUeuvAHhcWftRa26jUzreyKEaAeDd3
AFGH0M8K0dCMUyLJHeBsGBtLFOSlPqtGOGWDNWgSlJ6YZEjDqqJZQntwXXkfs1OCoFYvUp//dPGj
ie75JGG0V71BFDMS+HDo/1UPc7XJDPpSFpVgvi800yLN0b7vxraMyejjWcg5xFxX4T/pw4kg2dhd
XuxHtVrkDCTWY37rUtGMuJykp3h+8ItxvudCgUSg2S0etT+MJTxhJStAJaD+NFnmSJESnBySRgAj
cmhgUsmZRZHxXRsm8RRjYYoEIIHEQiieCY/Xq9VfFV3RJ+rRbzdhvHImE9GHkcbbpj3XfGiTNU7p
5Jcc4laYmvFtgl2+J/tCFDdWmddjUMbLKJid4SD66hYciL7wCLLrSfBAO4Z1icMWI7tvDDZ7FEuk
e2bdK9utWPpOJbt6jFcc1smu7LRT8yZjTYgoknc90OLLt1gqPn9PQUbO9bFGnia091eJzDkmT9Ts
bQQFajcRZetCkpLQ59fGpV+tsb+cKEqkMqgde7TNxVIXGofUp4Dx3DdmYzZ9SYfBF5M4BY9QfwBr
klcRexs7M4uVeVYiRZ2MAIzQxJQDz14uzVWIVuyn/BO60bBS5c+XqnGopQ6oh07NE3kVkDXETtnN
hl3OT6AuyvrQWf+LJQSbYpZInN5apUBQkLJ7QQgS187cRot1LeshcGdVvdgYqrkWV7WXlQ307V+m
EO4gL/V3axkevb6LpvO5lUDI73fSwVz+3UKwaGlFCJ9GxikNX75/EoKuZQaUiYZ/J5nnRvy07/GK
xpDlWrkoNXvQb/cqWEQRDDaTbqCZtJy338FbPVpbw5WDFXBScL3s8yfm9PVC1gjYhNsXj/eF+WQN
52TMV1NmGEh1LDl8+xFtR5wA+5kQpSSk35xaWwSjvvYINbyi2HxAf298T+HqUKqnKPKczBeBN4hI
/rcezMz4n1dU8VeqfVX2M5ph1rVM3Osc35IPYJFIlW9mJWdyVhPQjkqOb2CH0PFWA61X8VpoCkHc
t4/E78dylQ0VXMMCU+MFJy86d+ul+eppReg1AcuBMpkofkzY4ZtMG7weD3qmQdQ6bB7MoTTpoZLd
Ip3eHUEiR9ORpl3gdnfubsCfQKc7zMJHaJbmpjE3/gdd2luQ2WczQrOKwr44Zm+1DcWQWg33aA/q
GbNmDqfZHisZAMBtVFy3hf1q9hXCxiEPEbzkL1kS/i00zt2HUXDJV9LbmhaTfBr7HhnpjpStK86/
HqV0FWnwJceNYtndv4v9NUvWibCBytQ/4XlzQgigEpRpQ+fxvrQ0EM1hrKWjC2nsZ4KbigcwWkI0
xqKfRJsKvQoNNcaVE4aNsCIvRcWLqBlOu8iJMy56K8lUebc0sZ/bFLca31KE+aLvUKCV+42RG9A+
Uz91/7BqKwBSpIW9azILSe6P2GOU2vbyxWpehIKxeOIeWcQijR7S4xZ+Ti4KjzqumfeSSqGS9cXK
VgonTGxe1YOsdo7mCyjNF8YnrsQq5szewZ+ichS3KiJCU/TX5ufeIWsqmygHCjTMfTZXiSQ02hG/
upbupXXY7bq5wCgYAhgsnSH361s1hUsjdK8Bds4rkGwpeFf6bBrxgKsa6D+yVtWghXZoM/RJ6usq
q+rMg6NYYrmqXMrKn2IDZk2eTll8uN1q0dr9TdZsYx7SPQ6FvWwX35j2EreVm9orQQsN+3oJAyEc
L8htElUdoFN5RhqWTULjfwbU4x3NofU08gCZUZsp+Fsgu2mvmsU8/4f/OBECLph3uE6+FjW5vYtr
grUdP5zLw0IBJS0X5UHAqWavtVvYJKw3Rar0BIaRqKQgIiyLh1fcSzpsdVL4mB9+rfrSn9il+2p6
rQ/iEG7sOE4lRkotex98mdO4TZtnD0JJJaQTBuJ9X60V28YY86GBH7bWYs0f45UPNloLRWbP2UVB
4WlqjYbUnPKxyXdEFVo6rjd2iwTJt7LvcEah3AZPZYKFribx+PsvlEQzVsskYWCaS2qB/aOXsrz6
QgK/o2QCo8Lz1XhY3A1obakB7NmN2aPQDoHA70uU8njvkGFF7keN7VJQxPzu5niBdzs4DiKK7oRH
6+tK5QyV3JzlCRdvWs1BDh+0t2iZeL+mpN3cDi6IkUbGlk41WtrJ0T+lue4le/0o9Kpafiukb6wP
cRNIoaHWkM8c46+O8f2se69db2IKghbtODH8miaM9RrfH/IN7PQka3VVAxQXyq23IJrUrFDiOD8R
FdUutvgDLoWHLlwd0ZkI0TxU7Bw/YGhsXIs9ZHhEJCL8AgP8U3QXiXp7F0lFLGe2eDUlqHlfU5Gl
xNTXsKGs8TXY+7bnVzr0WJePxELRKlM44Tae/aMkXRCOSlacTEW+rdLWRYi2Ia0nnDFcLItQZdEx
77ZH85MYdjWei4cdgrrG4mgyDdaUXx2+sA7zLNFaoy52flq06+jexZEYMxl9Di8/5L9tavScnoj0
vvRkqs1Vh+7QoucAUNovaRGxmAaIypIAyOkOpFkLf4LtKh0HERzrFOzISHC/W9YZm//thWtAF60b
bWgQYCjFvz8l7h4mEexp40BgGr5otoaCNV9tVscTJjJKVtcfDrmlJeAAxgAPOvdqQ3swy5N3kUCi
GLJgm2NP+jE3YyDduYg68fvxdpclD7kvC9pTh9eQJkQ+C45dtMzKp3lUeAoZ5gSP1sm0qmNy7Et+
PvI2g9K47ygxJ4XLvjPQcMDZ8kQBUgOdgZ9GTAm0muviC3hIKxz2HNDrXFUh7PlvkCKOHTh70a/p
oIsU6yY5VuHEQwuLldXfPWEHciK1SGxm96/5j9WI9byhHhJlB/RCHrjmE8Oqw3fcpdspQ2lOwftR
6KSvQhb73GvfbRbshZykZdY6qktBrubacNfZiY9a8kwQGUWCZeZEQKmswaeiLL+oOg/nverRkj6g
qp/hQ1SXxPGq0RQX2VEveS8hDKVSzgGsP/DGa6xWmtXEteFch63NzIJZG9dJTLBW6SVH5+xs8dmr
zKoJQDt9svLZVtdJ2Oa5RyTDZjkauwD/9ZqB8G362nk8WeXli3Za0QjLOpumnTYap+pKW5VYS4rr
GWjma+OZ6cXkDSBjIMhJFXRUgHbSfoL8NfuP0qHMGDBFyHPCK9lafBEoQNUrmxPvVGM9/y4+Rndu
ng98VH4qrwDo93swWkmWw/0FGmuGQz9iOTPrM5mXSa5oEGRiXa4eKwLO2PQ0i439Hhr9hAHGEi6x
xxElISfiNNWmHwiopohm+zCcHfqK30wM4tt0RxzlGvwuQWhg3UlzpXOFuT8W2jqDiIvY4L5pPjmo
dWvzE29MD5f/dQB89MNI7tUASdVlxNnB0lzqwSd2rdpWnwMHeuP3EXF9MG6aMxJdNVI/6xEZchhD
/dPbZb2VjFu/OnEdGp7sn/e4NMb9EuW/B9EVu4kAQWvCvjRdwigfGsNn/M3ZQWyGnhDt1Cy63x/C
OqrBnQxGy95b5ZZXnlKpGqbnHVPSNIRumh0XRBRF8tBWV84rGjgPsyfgTfx2BwxIEgVUAhVwAg/d
4b+na2bmLhlcHbJgJ/NNpZ7GD2FnZY6qenIaPVgQf1Ru0YVC3DysLgkBfdSZPyzQBCAvY7kDaERp
SkIjHoFtH5GtYef5V/5TsLQWRugrahaaWIzYN1Km17m3q9ybt0V5suCTIy0uSWD2dzocJeTi7LGk
3LWqH5CdS8NIFNqxUp0GfOwEuETr6pUgHr2T8+YT+8ZRZxQKfNvPNWzsTESSiSbFMFkNUk9GJxSk
ZYjWsqiavSdre7fidtlMVoS5SQdcGJ776laPZcvyEp6hh991ulGRriRMIPNRqcge6gWb+OSjh3sz
MhUwPz4YuvFPXgkEerFMjUFnK42V0aA3bmFUuotCG+z+quL2JPPfGkQX44tFA2z148yUELJGH8/8
ksiMXyMDVBCQ5hfT5rakPwEcFrA9Tdq8vaGCVqsUKf7XxC4ckWnlQF7sjHq4FQDtpRsgG1y0zQWp
CQ/zmDTenrMOduv3RS4Umi+3vyLaz/1xjqWdthaWQRAqFuR++eqn1whhwEyq2UARNV5cnhCtbUwG
vLrxZnJCP8WMTBzvVXPBauVmZIMUO5goZObsZBACNw3AoCvmhTNmwZ16KE8fezf3ouig6aO/zVHK
YvHAp+pQ9PM0itrXze5gEZ1CRdY6RWuSdiL/Pn9oKQNxaLx+8MYquUNqRC7PZ+hs6gkEep3Fzp+g
Xn1BJpbTCiM3lBkO3a64AYiZfo0IsjRhYh9+b81NRrScI7HxuH7sNS7BJvYNPbw+A3q42TWL+pj2
c+19D/BQ4CcTLtYApr6JjV2bFkH1l7H9beRfc92EAK3IE4UHA/cwYJXuf+A/dFgJreIGnPo4+EJj
7+e/CATjE9Zfm6QQOvXKJQXl4peT+Nkr72qQKQtVHHaSXpivb5q/wSvJVlKY6WDMDAutuEIySJjB
tSEpmWjW/5NtMa5XC3vAe92FdatyothFeOtRBeCNIsmeXbgFRWh5QrVlHXQjTa1arNP1tUfzyLBc
aOmB4ZsWtWt/gpmENji7UTjIB9TwwjwUlW2TCSs6djizvffnGgdu0MsS4VYj5ridvvKMhXsT3TrS
dAz1/UoqiojbHX8u5NMekESbJ1zAjXP4KvlDQP+qDFu6awEo9XPtVf1SZD4x4psXeF5x0aCQVfmy
NNQGvgizMOpfXViSmX/iUxeed/7YYX/Hqd2fcDTbFAB33J4YMQcsruAM4wzwSZp3xjWaMPna46Ob
pJiVYZw+Un/4L7Uap32pUje7JZaDAE9MVicCCMsQPFtCJexVCaRkpXOk81cnSViICrS8rkjrGzCn
t9A3o0KxbMuixC79SIizj3YdsMEUgoMZm+O0+P1ePfvKO3x2DMoEytwEpu4N2Tmlte/u0GYB1OFk
v+ZoTdAkxD/x0F4PZ2H5pprx7xuT7KqlpRhcTECk/CfALOllW0gKbfBtprj8VnQjtGC1AwJrAwaQ
HQGb88xG17foftHyy2ZE96y0ERjYj9vA3eikMopdo6uo6KSRS+aYSYsLPyYyN8xmSOjn+4WocEXf
o5SmeEELjAFMj5l5v71+rIyQjU5iG0mAH94LNNjr9OlwKNs176jJ7Ua0ntA/+JKRj3zZPuUB0SjF
rYsWTzrczvRc9KaRb8jjyNRJ7vHGnkVQux+iWJqQdqXeFxwQ9ueLd9S8mWV5LDOpHPikxbb/Pp6O
Gztog3A7N9Z9HrmZ34y36wncJMOSNtIAYNEJFzLU3FKEyafhHwPY2GqC+pXI4RlLOX5eqtRv0tzB
7O5FmXutt9iYnpRGxJPOFLXm5YvC8749USqYO85cWp+y+x+SDteiYBoB0TCp31O3jAoQgOrxdOg5
COKHcw9zk0HVnxmXnGcnJNMD6klPLPJ32V/Ku1n7p7lKs3GGOi/V+9o1rb9HdABjfirg/5W5zvkm
F4OLdfcOTzqBjpw74GyBk4Ne90sY34kTf7QuJzVDelahWiAuYoEsqHysmNSDz6Urdx6sg5Oy9xTZ
iSiuDsc+JrGI6EoZEWqCLG1A1BADEOrVOD0hr5x9ltkkqnfc54xlStbAgxF2y6BCdbn33WkC4xIy
TtnugQ33SG4Pg6HIIsIYNf5szzAF6ETpTun0wnJ8E+wOMgR8++Xhu/E1r0kGL7UDLKhbWoRUHZjV
aF5CvlHrtOmyfrG8w66v2F00aPN0LDHQs2yRqsqmwZTi3z3OqHW2akuNUvD4sBbQBoc+iENrBlxW
FWuegGms466uKArexH++a+vDsc2uiew+dQf6kiNiJv15dPYVMC6OqT95aT7pjv+4wwKOYyRXRkeU
GN3xQaxBVNl8R460MgwhXUi68XXLElz5QkvqcUDpv3uOfNK+cZhTQY0CnLN3ASoemHQl8y5f4GKi
tkTqlo1X9lB4dlOdWJ0S2M+/zTvPZSicFXg5hP4Bzeuu+c0/ZjrxPb8b5MrclijpwnJ0R1TLvxV5
fX3fMnl5RYq+AFBEJTzqHgalFAf2QeCET668uGh88u+9Bo7iEnI6n/uSHIClLUt0y15u5+cTiwty
j7DDtsYqo4tyLDq3/tXcGUaGQM66FlG61aojyMgjN0pVSYNnjMMgLxqXun5gqcA0p2TLXFftX22S
lv7UN5PBxqSNyrsaj7uZrm//mSOw2Q3V4xFaPQ/ErbiuZm6zaRzDjeRpShJQcEpkiz4rTKgdcLf6
uha0NtQERJRCA8lRPWKF1T8Lfok346C3cZUmIhOqF70FFTD+iI0+8kDrLPyv+ZT/AGFiLWsBYbBF
yRDYSXVhmvmdCdAnWRPoar5VL2qRLwsuVxNMEtI2C8Gc27OedwrBJzUtIn+3gFNjm1fdoAXG7sXc
XEWsqgv7Q3Nfp3R8ESVdGLIjaDufr7dJhRPSpK6Nfs7N7tVoINxZpWrHbOCbdjTWFk21Z/U5VP9g
8R/jStgQkIz2PNCCJVppkRU3+aTNN+f2Nmx5vdevREg4MyUBINtYEY1MdcCwARO7Vubapm6IPqjK
bi2dk43vyGh9dGfANEHPkZR2Xpz2aZdqKJVBLeRxOlkC17ZHBqNBdWRdI48ZogtH/9mDr7qlXcfo
kRoRGjT6JjjbyGKuHOZzVJm81D6nIscPllPophdwT1ED9WFlOXnTBHpVhI2s2Xtcb053dEpuuoOo
XFYTo00tCyyhR+qhoJoV0GNQdjnmVR1p/U8PCycbQu1GUaIreW5WBPm0XKF0tPKaAPqrAxjFNggr
DTAoPTREUeNYBkFb1ps5dRyqQhOJILONazuHpx2ppOt8A03aObfrrEfLiDYcSM9ags2EChvYlpd5
qZL7fjeD88yxKiEQznXwOJZUwIN+tcx5v0Jmix44aTBZ0o7W8LfmKzEWv/urTlbAnjYwo6ZybkSP
54JebLXlRRPhp5zLax8DPhWG+K+Go6hGZFnuIeEGGqr2eXdIS7e7gFdRBW+GeYCPWNJNLRGguWM9
Ch0baIKLTsXoC0Mwh0ZTN/ptmVCWYUvgBVzgz0dGC16VSZkO2gAr2mCqRaXCunLlV8oEXhwxsk/5
w89oLE8oV7tflbt/o4JD0yebrdOWbe/M0HgoPI1F5+HEMh83lGhzuG/BPwcit2No4os6BNCRWjOM
FY/yj5R5fZI2lACodhT7vOK1UUw15nrFrncVNgS7NK+c/HTuiQ6UECIYgcg12+HYqa57EwpHIvr/
/BDjdiiKd3LaiHUDas+JXm7IMPfSQ+RQ/uT0mNOrxLCgO8R0dZ51eTbeX7Frv8Ggg3aSzUOq3c0z
4rxrDqjwHZLzLUPBGllEw3IWyU1XB//zt/+AGjcAC+lyfxk3EXNyhhz/C9W+f+lossn3mxaaXM9J
lnERi2sixLH5VZDlwvWmyb4o87YffzhMQ7hHm4WOIH/JSOyLYB4xi54UzNtaOK8+h6TsyJIIZyX7
rq3nTDgJMza3XRy9JdSbbM9/Qv0pVtwFE6w6eMXfNYSjEFIeTyL+D/CkpaTwUTncu/cUT5nPSaH4
vzXTu8kfNQJlSfJ3lTr9o2JzKujAB4wCGu/1LHBb8SGy49lnfZVWmZKBfw2Fpt1NBqPVnH3c1pxA
w4JjIcUY0k4efl4MPr9AnIpl9EaBPsmyeG9JeEhqCjJXO934NySQxQwvUJRdVYxZ075zPplKbjLD
rOrZXaQ7LhHC85fPIL/saTENEHo/bfFZ/5Qvn89TVe8prtdU36o1zpf2nz1XpnykvzoKy2UuUYDU
igQaRPLGGhWEwVm1r3x9Uu/3EPzDwK1dzN9N39HBXwLa91Y66VBP5zsv1Ox/fvVxtyC351Ehfd98
SmEFqRQ1ZLbdcSg6oBlkFQR2uMC2/8awBKziwJNmYHT4I1ZgnqXQrfHFES951akTmS9L9YfOm17A
nL+4RiOFUrKTdYBTDKl9PtoiGnsIncCTeNdrLG/kDclPTI55ZQhArUopp+D+/dfVyDH7kcepBcBC
bbxSutiYZmsHBYV6DNeLwWDeHOJUSHFNcDz+q7ABT+HypY86wWrTHxl2ru+IcxfjT7qhWTp7LFU4
ucjdswQgvFOj5KXUsishQ1Ayx/gMjyIj7bXwjRuKavIlk1Y1taVW3X5599ZSUB/YmaIRKXmJYr4E
dxXbQOVSRC7oE4cjw+D4GB+tjbzCQSMbmxEP9s36U6lo7kbGMg/qUuP7qoHCOg2j3W28p+Ejhaxi
3W4rUv3ouZjSALobAEJWxO9LF92exxW9quKK7KyAobBo07KVI6CdZrmE2OwPwC7kd0NDItVVCrdU
jSTstVJoheSQUr87+bvRVoey87J30uNnRTABF5ipVm4G40FdI2brkiBf8ZuycAwLQzW/f9ob+v1z
g15MZseJAw5wVHvqoVuLQSCwPmWjM1vuzTLSslcw6sSgSewIXURcxXXhHP/Sj2VvqPeEuMiCaLg+
zo4KUyds00+M+iTaVBXYjQO6lCnTZo29EK0V/2aQuQOmNc5a7barA40UmY8+T0gKf9PmZhlPS1Ix
tqSkkOBfCjytmWHcWKWB+oqV+3bZ6F8acTtNIKusFCv9IaY1K7jpQAW+VAt+MJlu0+vSHAPy+qtJ
usN7b/8CIVZSRIkBW5RIlwalgtUoPJgu6jGCdw//T/sVwk6dbkGWFpcgjePMAyNnrMAiK3OeX91r
Fz67OYqnArP9PEs10lTpiD/Wne13zn0bf2UMkM7YI2llKGevGYVtCyUoIlx6bmWLA1rB0BJ3QUtq
BrwH96xCtU3awdxBL8L2aNzAEhqICE3eLS5JpmE6uEYqTf866HkfMdqpVrT8Bey/M+f7FO15tkcH
d7dJNrFGHiHmzu5PqBAQaGZzzkj35+ioyMegwPWFWfqS2FDFsBPvdS+3E4o9FDOfWYSzISSiJdrt
ujgpmD1YgyfdI4wr8dSn875g3uXuI6U7UQH6gTu6l+649Ana+9RiNQTLIcguqysoYKJD2p98Iu8u
5ukzecn/RhVo/8ysdr7m6VqHgaVY2lq25kNDbG50DvtJzwylL5AT+xu6MpyF++tpERSHsX8HOtbf
wxSQnD7J11VyOZlbp63olVQXSkDP8jWt/43NegiCetlExThzCr7AMbTBTXkO1Z1gG+1C0i/6lMsb
9HFADL89Sjaaqc57/PZDLO7w+M3FflDO2waUp2UXOA4uFFv2ih63LnsPNwJAg5ROv9EaHf5NzOUD
npAFraQs0KbOwLSui7/WJ7amuVw/dOOD0a8mBD6Sg9QTaAhbsDPU3vkk2dYuSKBANJ6fLwwqh/Is
iaSQuWHNKxIv0sDsatTI6XLODB1vk1edk/gOBc1ndcu4JriEzWxwzSdUsuhwgYX6gy4hh94lWxIu
ToHZsIG5aUC6Ll3PnvZUqBZQ22Qzm1ND75AwVD9M81doh1aSbRh8EyO15kpMGixYE9R4dLqWSHDV
40Pf6MDTNyelB/YBnr+gZkdAVyI8ilSROZwErfSRn/OdxGLhNMmpU2R4SCq/AM+Nqwp49eZScxg1
fe04rFTBpcYMkdy+BsFLAFQzPpuNcUUJuAd/mmY6BWp1pxGvLNGLOfYIIsxQ9Ebzc37iaWrL/ZIn
LY7Jk5h25dU7CGK3shT4hb5c5uh13POqv4MPmhdMKQjENXKZuK3mgFWL6AbIpVHvX9jopucRsl86
Ba5r/IHW8jp3I5/Q8wQU51uQ3qyfoesqSjaoOTUjXRSWo3DjOu5L+MZZgPpoHweOudAh9W49G5u+
Q8Rd7fwlY9O6pbleQFFG0ceBuk2MORdLVRjZOHXfriDK0zRCwfm4LzxJXyOM8YHDyKBx+dq8M6Vr
5JO3nerf7xw+luMMrJt3nfCEWhxlJ4DTdJmo4QWYMc3vsJ5XUpD/IGKvxsS02TQWHa7uiUsxCKaf
H7qEL2jUYw9IBdrxM2YyYdkV5+COJ9Ovs6ST0uGHE3KXXHWnEolJ/nyAMEOmDmnxgas7bshG3hZS
X197o782m0Sx5UxRZX8rN8AG5sDPFg7401jRU2kLu9C/VdS3BVEN2W+FfHZz8/TziFe+6hm0Y5C5
H3s/DgXk2MMrnicnIROfF/YyT/aYNMsY3cOuHNZUEnZsfnWsF8OJwrx/2Jpx4f5NT/NwBC9C6a9x
OhXv+wpoxmusRjwXHeZPltiFySYr6/7PWZXxuvDFOCQ1k/1qkSgIXrFD3K6IWTU/Ibpoy4gH4F+/
j5tEA4tpcEXf/Rtg2L/tstXPDO/V9nDo6ICLGNEw8RmCXfS9moxsOkLzY2eipC47JKImpcdoUHqD
bvYZEnGoRk3jxPmMsg4R3p6ljSRosUbwcRR1fI1j7IjYv7lgD1DM7/bwC4jCkp8tX+qtghF2Mc1r
V9gNz6NO16pm4p7G9drRZLY9jY4Lg5vUe9zhzjhGElNtwH8DBV1oyBXXLzvrWsuHkJ/dgZZUUKzn
oDkp0ZRckGJd6ixwsvyQ9pzb4rud4lIqQs7X9dJ2U5r+EfwVoKTLq5zJFc79embPihlwEAqU+XUJ
BWGGFXDN817KuN9MiDHBftbr2LLVzQh0YMWP6LI2FZUgNmOgZtnxXbNGrse7GP301fJ1GOnKjqJC
s+PPrH9WRj4ZhFTtV1Vmjk+FURutfuO0ww0OgoCfISMVZSjYdGGMG9mmVe+0T3BANc8szMYhNMPv
Ht1xNTTa4IX/lVr23XB+qYtcz9KxiJZ24VTGrBvWQelNt37CI7hROc6WmQnKGtwsY/ORIZ3pIycB
8RUv2MhtKak6tGv+e4Sxs3qPZGgH+JLVAwC/1VNHvkHszfoAXe3orlo96J//uwdxi6ROvxDGCbQb
YXvYOVnaY9mUSxYzHokJaYmTFkNOF7Aou4vKKwakGqVVyBcUnwqxYQ2gXi9Rok2nQRyqNEx6QMEU
UUnDnSma9pv+mJ6LL6f1/HzeLYKWw36rKUYKKKQ2kyzn4Fo0Ui6yrjG1jBasLWB1mQnNoqlSn/89
luHLTGzZf8AuiXZ28Y/uikqr1xpnd6bEllNLPTTbs/tirmln5sAuMX5/exACUVisVydPJ5T/Oe9o
p5uvYIHIi2ZPBb6BZhxmgFwhkYCA1H+Gvgz8TkapthZbklm8NYD5lSIE2SyKKy1OTCCtw82u2NJh
oxEcdjqgVusPmI2kfZjGfwzJgDbB6YoQNF58i2xG4ZiYCg0guiaHz8pvaxW5R4+qK75lX/gYoft8
Xda7efobB7nZgUXhkG7+GGNlcXvyDgASGXLKwiwFyz0PTkaF44yIN2h+aQ2alkEQcDNIkNaS81Nl
+j883ePOvLvPx5LIIZwOH1mFvkf21WcsHsDYcL8nXAiN6SdB98L4xNo47RpiOUIgjZhvxdyLSJ9M
K3HSB+HVZfa3LN8M74Se5AE/lIN9EV8gXxaHQOUGh5w0Q9njjDTEAd2EOeGLNzmtCS8aGPQ+WFAe
3QRc2L23dDPRuzfPfvS/25R7ne4Z4KIW+kcBA7qcB5KY8+n77GlJ2jZnOntnaotetXOu4RfzHVzk
TNTcQQ0PcVKUfJdn9GR+Baw2UqGu3iPQdrFtNXUoy+iklJZGsBVg554ny5dYZUZngVxKhf5GzRIA
ypLVgPggxtjilQIeJqjy/zHGE6GWuNH/3zLnn3RCWH7kv38Bf7EZYPKMemW0q9QeNTL5UASw3aIM
4ez1rOwAYqe9qaFfRfy6C+cATa3P2JhUqyiHiG6PIo/A6cu9yFNAG5r0NHFVKT+YsxsNA4ORHJ4q
XNCDHDEmDhQT1RjWxdnSo0pAJfmsIgzqVzIKpZUyA72Wwm4B47DZYoUi5P1iFHpU7EcGfiELPKQ6
5K2NrZ6505oh8y718MGGjxYuW9hZI/vUrz6C2XqNRtfXoGkV50okvEozdLEF4GPqdppg5W94Bwd1
OwaP5mPMP1FR50viFTmA6rl75Dp6Vp5UcVQk45+xl+Nu/5ikS/paUnwO2Dbgt5bQDd87C5sJogTJ
DZxm+9UmcJh9wJ1uufmb15XJe8FQu4wV3UvG1yAAruOXkDV5jwMPwe6MNACVpTyZxHWNKJBDve3s
MA0Dhsclxf2qlR979W/ZmCRZIVbsrM78EHfo82blSHInIqzp38ryBhwPvbCcoOieMdSLOye7CETI
ZXrqeW2GpSWz8T5iwfcRkvmIuH/INrD3oPkrExv1ShM5xcHZjo5cg4Y+lB9Y+O46viruI32mpvjG
SYAENv+Qz3G4o0znJgXVfYyfcrtAN6yDz7KXy6dS0chojUc7xagbDC5Ee0bJH0U7YexfM95aMzVL
L2GQH6u6Ea+yArt+RkpJbt7ldgXXlViaw0hPpFaL+RkouAOsarJpkxPqAgxmec90e5xjYNYPDd1C
Gk6d6KAauMzDZ0cHli+sCLQeTw7nG4qgVjL7SNiRLWsueBxYq0tvRLsAf46jai8wvlOp7xYM8T+i
ydEHN14KtgWhQbfDeAqtJplNWjnGuIOjFf+YL5Mxa327XnS7UJ0jVr8VgXIHfrXvUwREPEgZcWYU
6/69gpWbdFdq0Lbvrtzk7+Lr5HTZTTROVmaAqwfdV0w5W2LAorSicLac0iPRF3uexBtW88jZFQ9w
Fol4Wo0f88MNW1ugXRM+bh4xxLPIgVhcOIwHUdSLumOhc7n+m0DzcP7Wr6BvJd35mwW+oFh26+84
gUdX3v/AW6WHkMWH0cfOxHqhIWl+4iYBUvxZbK6Mj5zMSnsgp7Sw/aVWY2igafZmuebdClN0zFj2
7QwX4wAksDqi6BGulArbaulqTyWJfe2EaRIk1zlKk5SZigCDf6Ftg6qxUOy3Qinaqh2uPr40LcQL
zHD347IOb+piqYnGEua0SmNP+L7G6YTO6a9SqLf9uHunRp/kiE27QreSVV0MnfdHSN04AzQUW1Xi
3kZ/KHij2d1Gi+VhZRZo7hwLYwi2ZestZsCBgx1/964f7hALMe4d+Pbm7H5wGBMZLNZvsRl3T2ng
OHwBiBI0PMol8U3fOv//tW83H80FDmuo7Jq35U0+laoSqb7rnn6AZoOh/U1d7CgSVnlS5XfrDhpV
dWWa6DEXY/2LWCxL7CCK2FHxD9TywYVHCoX2Pmx9EO/qITPBsjBP9CK32SJVLWsOoZfHE0e62tS8
224D3UjXJLM5plQpcvFYftEa60g4FUDuJX/s7PpjKDyJSQnDpBgc9/Ldo+Z/i7CzFpHG9QLemnzP
AgZsEHYfoTDPD5UJpFHeccbcfwVJgThvPIciVLzBuGzlIz9CnfAhRTWyjrFyBCDk3TyKgbUCNaJV
zpy1wT1DzrwNf4pOnz+iIUYOQvA7NZAQfSa+aViqb5/aDb5y3P2GHeb3WyK+cxceBXHIWomDlPvC
NsDxM0LNx0cfqnqDIaEW7oxzB4MfV4uBI4vuYtaJe6yuDrLTW7gr7YNpIXuyupyLRVdNFKxTzHtx
hoTpxQk03K6KH6rruyQmk7fgG4oJNbpu/D9y08zVk6Fr0AczOyrjAOGwz0HzvdxWcF/EcvholSui
fcmGO0m0cGarhttEkq2aWIvr4s/Lk72P3t/603FfOo2U5uBUVvrTaxIkyMyCepDgt0V/GJzbeZn2
haJW3iXISzhwf2RmdXKFpAc9cx9CkhJ5ZVPXQkSFSzTSiQ6G88M4lhPQRPTLaAJPA/3vcBhaSOho
4dFC8+IGlnaR30i1UrLB1PJ0JK/xNadaD+uOnKDLon30nifrnf89JJZzoYYN5+jKVEW4Iisebres
wTpVgjJy1E+FHPZzzSLVh1bTgxty0qSP+YEQ5LywUpx2XpR0Y5a1MR92XvDg3DbRM1dgjHm2nBc1
YeQSfI2itU2AHZuICordjlfLXmTnXpTqS6aJIj2/EfXz+KqZ5VFEIxLKkHtTeTavxHdaAInAwTUk
5Ay7FYhZlq6WkYEJCNhbRiiVjY3JwNhT6pQuWr+ic93QqFfzblvL/4i3vDZHorXokdbssBuuk5cV
Th5ysH0rNFCe+1HsTDQ7jzGbZl6EM7jso1TILtgq8TzDDn1sz4mc7AzNn8CBnLmnbQa7Q64cZX2d
9X9GkuYMR0OcSxWnmFATFevfLXn0VL2RTroph4FUPgjOl4K+NF81EBUQIA7Hs8aoEz4IRuMFsmmp
8ozzCmH6z30u8ere1xUncOyWIsRxHWkKlKSwnzAwxXBAzoQeuImf+SdlKaCsqLLfqLeuSzdstUqS
A9SpOi4S6oDwHrwAppFg7PYQes7JtdXYsyKmAJCbg1ZTwCPhjUDHbZg0mA6yBB0cWEg76okzeaw2
aTSrv/2suUjT/tNjMSIVYSZmkA7iL/xOnh6lteICo03IDptkLnaHIMHfzDSyYf08iZDdaBRkQ/ph
+pukKOIO/YQe683P9cJu+87EdaSfgqh6+a6XJ6AVh98Y2t9wkh2hQa2T/AEBApK8Sz29SVvLjsAU
vvurGkG0SrUEhlpy2urJv53Svh5fib3nh1bOnzXf3TMLy1mhaOwlE2Cur5o7FUFpEVlag0vJIp3/
oUP37UjqsvTHnJ/6RoG/a4vZuTN5tbkoqUp0R6JClp6x+z+dnO0on9HDhPpi7LL7zjMZVXQWcfEQ
1ROOwPCDiQkCyg6XeMkkD0qC0xjX40OqT2sLnpNv/ZbEbPOIR6T+B1bHvNHPFExxQXDMt7vkfWvA
VTfkc5mM3Vpq6trx61DjlyDyT6dlIFHmlCkjtrvLCMefaQ253nfAGtxC9ilkA21Kb537YdLKQEXa
ID8IWH0uKfzQDLg3dTolY/tgp2SSKj87b7V3Z6IphTbJj/9sziQNDnfU2YLRTp6bp6okB2cuajtu
zZlyGCnTBiFdfJeb0qh2BfgpVukQWb5etx8pRhuHlCEfUCdlXiPleYgw0/jDV+d8/0AP0HghvZ9+
bAPREFpdlk00Q4P7Hcg10estZ7nu6eHR+krb3z1kybT19ohmkjynU3u3p9ELhSyoXswyIToo2ybn
+czTpR3fM1TtOzeBS3c41RQr6GfSqCtKU+a2Bk6wKpDCsJFXGIN4tNGxsC9sdJdJUEFdyzMhYrF4
S8Y1A3h7Sxeo72Qq/Gg07MkWzDo16FqUv6BKwCKkUHRXpJQEUcdAnhlh0cZpF7L2ObUduvnGLnIB
mdQOxIOGvLSTKevRbnmbv3PCTLrgtFvFk5CWSH9X97iTMWv68YDOsivvKjKenmjgPs6U4P6WWNAs
2zHoV4BKcisPbAloLMCkkLCvBi5E6/syb5TBQDri9knTZxdzmeg6D1YYs4eVFr/HZHBJs81j6JeP
ogmhT66W1jekgZngCpwP1EE3YfrvvkGmqyEYxmXPV+2VJsdNGfPYaY415uHmG+wJG4WtcHZQ1sdb
uYep/OxAehoek4cOniAs0/RleJ+C4gapbSh3X7AT8j4Apss0fJNIbi++9EXhOX7eGukQDAiCAD5Y
vLDsulONEmWgVv5rgLyDLVIG/UNk6ig1uM1x/zZEWNhW/FZo09dpxX3hSqzdXpkNjpGkFGX1AqOD
MReEBtUVDRQWFmOZQ/HEVnnyw/pcDormx/Db2jXY3uRs4g8q21rvgmh8M6ZPeyOlq+ofhDIB3gU2
fnF+96Qw9kCnAJjTSaBOgLEeHQu+l8gMatrUaUPBkgFxcJPc4Ym6YxLkehkTANcJeZRdH1K+ylZ5
KKRUx6vRyjZ6KH19ZfSi1LUXTdXZCysIBw7VCfwWvHemV6Fue04xh3evsiP+C6hM3RxZ0UAct1uN
OlvwibtKHlp4OvfMXTFFgONd7Fs/Nlx5cRGwqGkWorVNHDJUuthrR8pJLShr5iFQAAav4JRKNXna
tV1cSwu8bera7VODq8mw5B0nd6sekwZaKORf9DaM1m02d5VvmgjXe5D8uGS8Bkb7ASPutg/s1Sw9
6OnkS3bUCxNQeoER0l8szUzE/zhRLKvHv1BaYlWUIXYMF3Sy9GK5tbCBPV3eIOVVv4sM/VU5pops
VzV7ZFhZ/2EWQXL1Y/sEQFSKk9FUu7IZk5hIJJtyFTVHk0L5j+JC9gFO3QRbSZ0LI4leqC6jx9v9
TWiuLbAKDW5g94BDPs5ASWdNhmYH0p8Vpn+p0On7v57dodJleqmDd5o/xejy9ae4hBs94QnUlkKd
5WgZCK09FLYohVsqhbsWGbAdnXqopPIlNVvWGBnlrIhlVg4Z+9gkTadxdHlCWFhOQVNC5isjucYn
hJkLBjpP9FNJZZPij/H6Nc/eKZcE9Vli2ddyK5lYU0w0MhsXBMhNWqyuy819gGXTycrHGGAZ2Yqx
HuN3yR4BmzsiTnpSsJGKqcG6tAcy0DGP962bgq6V860u7tr508mIxV3P6JyPsVSdE/8uPx6WVWr1
vVjB6IEnN2erhIlLvTLTDF7UXcOaH2Uh8mIXoAjdjZxzjLzLDRMlpXOypRCREB+0ucx0CrMnDA8y
rOxOskwf8pccr1u+1Z3TR0QOv492aquvaEswdewTpfCHeVTU+F2e3Rex1SMchTeJXxOsBELkq01v
3oxB1No48wU7+k1xz19Ite9+yx1plqnzdaknNg7JmHmqnfL/G0N52O38Z+GavtIyLXn9TuGJ8Ac1
5Lwalh57kYlDsgSiTa5p35iGi5ZBUuS4fYpzlTRnoxazs/qleun/sb1TqKR4rmQsdeKd1l+7asFk
8CDi4Z+H4MyclMoMI6zMnAKKmAO7FfaZpZtEEXTrtj/WbKKIJWFLXzghsBWZStR8Wi+U4XN4WUZ0
hnIdeREwyMdRzMNw2Uhv4InOvIalULTM64feUkCV1GG2qF81WHGaZeEc3TgOUVySlN3US2b8qtDs
SqWn0j0TLEp+3909CVsdqyiKQW947ZhoaTGqBftoKv7qGi29u8b9JvbZgsgxt1nsu6GtIJ4Pzvp0
IdPHYInQAwo0Y0H/WP1mbSNWIqA+yMSmWGgJoTZNT/fUYmhicB4u8VqeHqVIJ4NmGBgk47mc5P/d
kVRYkkePu12LsD4Kiap6SkCfUBBlNiLitAJZN5YFQ3Q9pCQIKiO0rWd3WaRKqslZ8Eap+pEBjJHR
VCfUkI3HRe2Eq6otdtCF8jsUB3qbHTHSuS6SSv4xE3hJ1g9qolYMI3D3x4iIht6OHoqhn77oV5jn
yGn2O2tw1vUMA45ZsaI141JL9nns8tkQcsA5OSDNU4TC0YfqJt2zpjRjUHIpxFjCFEgisso9Dn+2
fyv5tJ6rwwxflhcoM/+TXLE/io0PgQit7r0Yxh+6pJzwRYNS7xhyeZbEYYchPFFRaw7ycQu9D3B0
rJzEIr/3vdX2KY4Dq/XoD93/y8wIHskAw/ZJPiA8Fs3aw8xoeN8FCo/dmFF4ks+FpNGxtQJlbh+c
k3E1U3ffVcJKic7yd7v2bm0SrkxR+tmpFJv9QP6ixF5v5Vj/+0bO+MWlX4+BTiGA1qCc6UjhzyEy
gvE0EuyhlfhJxH6j+Yr+L+6vFyqnjz9zzQOIvn5OYn30u7cpxpwZImUFFjTQcInX/iF7zBtsKAN3
r+4OLfYJg35U/2pTo9+xl82e1r769OID0NGviF1gbL7FE/p0nlhNZlZS7YQTTaqTmJp9lmp3JK9M
UjMMDh/mrqamz95AFntYN1jnigqi3M2+DtDVHKFUsCyLDRUXimOn6F3FBl8GbBt/w6EL6cy2QO5O
iYLM3/jxUVtrEySIvQTY5QSxhia8E7+nE5S71tlfZ4CrFHBhmTVLCy+MxdZtAEQYk490HXKA4iyG
hETF4S3yRVsxgCHLg9xWVp7tIUsscwpz1/Djbl7EyuRLU1zlVCiPoWHVRQlKCSKRafe1WFx6kh8Q
A/iY3Sbz9dGlZ2WRf4hpQ7Z5TLI2lrmZxNAVZR6JyGLDyGcYonMSDwsJnT24EnNuSxQrWPbMyBvV
yEONtcSpxvZcr9ETfri4E/gyhlLseDjK070doEk/0Q+B+swFCZt4wQ7nsWJZxyeu9oRKzsEzYM1l
eQdEOrGQBo3yJ4EtsNPIWEBr1KKNLGhIkuz/C2WWbimvIT4suagB1CfrPjbB1jeQK3DSeZke6O0C
vdm95sY25fNz00DlxVWSFKHWleWIZ8q0oelfYXHfkeDVdtvgDhIUCkORTLfETBA2H52tAP9J4bgW
SfgHUwLYEdks9ZTzTVGgmm+iPbv4qOESOaWYJHE2KJeRw5nDmS+vhM0yDj1EMZzJhOn/JH4V81um
ldYYR0y2mqdTEJ+jEabX85wq+mURtVpscAPWL3N683rBiTkPlkMBTH8063bFO59A006zTjL8T15i
M6vJxxleYpj9NLJylXi9nM+a2M+UbqrDPeiHBdE0vuCOrPqfjS3wQHQ89KyNunpymiX3DpW2niWu
ZD5LoW2hwle7eg3aSsZEhfbQqzdJENb/iOeYixCuilnDdlaxM2rqscuIYpnGVFA0nsxTIGGDGgsJ
6POMkmPj8Zt7Mig/gQigu1HwJ1QLLf7ij5jWm5TgAK9XxrvECKKIkeCfIpggYB1Jb1Kw4sNs03Bs
0Psk8qDTMgfl8MZX5HvEMOXeczJPkK35joG2exlxiUsRYA1kJ7gCs+dysbC6Cu28NLHltmNRQMwO
NTUQGAHKy4abMOJTGvJmaNtOE1MY4v86WrlJ9AL7EfabLNP1fTNyLBvRzXV/YlJJTVinct8HZd58
NB+zTgkvCR+emVsmFHH53wGBE1ST0a5hAvcyxEMUQuYVCldK/G9m05OnvgWWEu2KDt30wzk896Gf
grNyxg0dRn50Xn5SfGT54V/Ki0rus6LS4xaGI4MA/ZO4zL3kEFGdw3x8yK3yVA7dfz/0sJrqXFAa
eu++5FtwyfDCyQr7G4BZmy20x7olFNoeACg6tb6hQTz2fhRG58JGp8WAI/63b+at4JAocdDreA24
U+KbJg4/Y19sIkYWh3Dy4AW9LWL0Zm/bVEIw9O9x9jAOGSjXoo5um7HbVEw/T/T3DWSHA7aYCsu6
TuC6STxjdJjqjXbWRYszdSnDiUZd+PFM3m3/HtQ4D5+ktZJQMGsGl6URUhKM04zSoFok1Rh4vUKV
Qbd5u0WO9rqfupjfiOpMjEEzyFlWwDIv3omjhMWhHra1dy/IPp5lrHx6axVJWSBJKT1/6aPx+7M/
kGTeRlmJ/cwZ/nXEvyjvAvgrrxmW83BTvsby6EU6826cmaqHir9HneQXBQdxJtD6g5ALP5rQRkk0
zvm6UkSdVq/RQMyESXKuYbp7tXPUdokzakoa25o/iU34yK4XzI17eXsETFnNGnwyEk+bmr8cVBgi
vESl0nA1OvuwQGbOa/Vx0itjQ6giL33ZhpOap4uFB+fzuwjnkkHoj9Kgc20okfqVHME/3fQcOiQE
X4LZRvCVopHQ0Uy1829SwzZDnSYlla3FXqKj/FTnNWgpr2rqTVZqkHPJj8nPaO0jCge6bDpyWlpZ
f4h7JZo9Ilo1f2kynjzPMT5Dul1C13KryERULuY2Fgy4fChtjRTyMW8nP6hbzA==
`protect end_protected
