-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kTFT8oTd85JA0I10fTqtZ8R4FV+GdXI18IQef4lG3Cr9vF1yOTRU4C9EG5em2hiBFjyQqudW2dsZ
xl1kCLbYgB4bissuKJ8WJ02RFlx02TyE3g4NQDqPWRfWfeJngpIYfvI6RpvPjFbvTybRV23R7/Yh
oMJGx975+N8gdaHQ2vznTknSa8bGZYErGzhq7TGq1nrVh1CDZ3oWCSAHdeV9VZs+QiMR9RLkroGN
Vuvz9EpqYVvzwmSmKTtPJvUgGgUOXkhbWwTG1ocwFSEbqD1IfMM15xqUv2vwVL+Tpf5DVSRFwpOm
2MDSAhddxVu5Hb+xFTf8Xp3Dn6a42jYrjShIoA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9760)
`protect data_block
CxEF4geE9HKU9/6pf4pUPmSMclVWmhheO7kb8eJ8TmOAO9TQ/vSsZs1XVF0k98WXqphN5LkeKsAs
r1AHO0EMAPhJiepHFsjaGcgxgA27E9r7UROHklC60LZK+2rWkqA1DdEdcu+JGKzHc1LOq71G77Xg
j8F7+ovKrzBrgoguPKjgq2pVuNWrEgAjB6KBnJmmb57kpIAJk1dvTGwYDzs6TyM6qAc3k1e+z+aH
2rAg1cyOtFKvoMPddsj9/kJD70HsT5Lss8n0tI39psK+V9GniqLW4XOE3ytu/j25ai5sblWiA+mP
PZr5tTOF5fl+0Z0aOtUU0O2CKHHMp2kVHUmA2JTqbts/qYor8g2qoxo1lBzlUoqSGhn6Oeb+kAZP
oH4xJHFJd7GTQTei0g+cLKIp5fQFO0W+p2SeG3iYJCPMO5NGX0wHJiZ5ot+3l99qIESojf31yjHL
YVUmw3jU+K32aWKF2h3DyKdxXE4f1th+HbpmwaRW1pDsAj1FmhP2cuk6Zqwi9Wf2hOUqSLpUSE2O
TMbR4wNxp5k9t5GOhcV3qISPchHUuFsqjjxAz9IS+zZliWvGncBO97OAlVh68o/lR7mNWukCP4eE
liL7TrSpjiuCsT0y1nvYWm0jIMID299JTM90gcIph8hXNkGRs2stDKh4XiNg6xBCiiqctMI6WWP+
kgKGlzNZKlFAIjqmLnDBLi+6Nu0f6U4hgOIba7qxqTbPCnboEkNFsZMMWsAuQB1bIMXh8y9Pb1FW
p4LbiiQg+Vhf/vfQyzZNCGEuguNNc7zaKbF7kJRG7lUA9GhrShOEBTWA07Ymjyj1nTA6obHW0c1R
eepAtc/MI6n1iH/Z3qRrJUMtxKairR4jVUOh+1Fuzhydl1Pbx8lWgrPX4w2Cq2jXIoEYCrW51uk3
5k8suKcdO1L/xSJJ18tnwGfPtPLchr0RrVb/GEDur1ZTwzUu90Yc6IRKHJ4QpaqljkYrdha/rBH9
3auqhOB0RZpqUbJADe1F2NJRUS0EV/MOxdfz1ATxJ1+Ahwh558P/1hR+HaZ5DeOL6IKIVfor+Y+C
vN8uj+CKIMzA7r1M51MS1mlNQLhrbWdrclQs3cy09B/HCQy8doKk8e7O0+vCpnfznAa+FG8421tk
etGm8AEL40UIZ+9fZpygpVVSCYAXNqL+HYJqsRCRBzml5zsuqb8kIL8d8gEK7xm4PjJ9I5nHqgsX
s4VD41d3ATmPRkm9XntRRiA9SXl7c9TDRuUsiCXjFjnNCwdYGSByDylk+GYjxMOI6SJMVHAvd5aL
FGSR87gWMGUpCyLuY5xRvYcScX0fODqwn6jRSvKCw6P/sN9XF2nfMs0uDjRAtg68ac1Ufq8BBgg3
/XZ3wYD2oOMFY+uDhiUzsySKKmt4pEycIPiOhOHMWx4d/HCoIPmTbmONIiwUkZ89d78IM+PJZ4xw
adD5x8Ep8MRl6p3PJBe2fTFmi0U98Y63yj+8CFMNxWVoY5tBzDb75/20ZwkNqU9aGZI6/wvCjzPd
tFxVKbwRbzPnw0aZrSCDrywigXr7STYI8G+iwQOfw0o1QBW7InUWBJEddlnIVUVCe+BYjq3wV6HY
oTkSG2eNAGzX7lQ9zynnGSxIUHoGctEJ/2INid5/ur2lBFGFT1LPRx3FSAoaCvBhL4BTPqAF6lr+
C4ChxcrdgB2XZ5jMBV7Ila7MgTfCMxexTLP6nOmwhW/47t6KwUVttS7Ek07UsvYSblaLzqxmH9m7
vDRUXsNywFnlBiNQRqa3JVW8yBgVquVvdN0GeksK1NEJjWR/e756D1idwboPzW4tym5Y9nG+krNT
xZSkme/KwDam1MhAS4BS9GbT50UykiwJ+XHS2/Ub/jZBYuDbLUIwflREp1qPcdQ8a7e5wGwZ/c6Y
mgbbKVqdsg+MsBzygZV8qTGiZPQ85HRE1f1mm+WQhaaZTg2t5I+7UL8buvtOxGAIUKTC4pcljuBY
5tomTWvR2d0zVEu/uX+kXWboZnM3f84EOPsJcmaSJMGCAH3rdYl9/SCBVg8fdMx634IJwKKEnxRr
FCguK1O4+C67Z5o70L7UQlp1d+WsHhxlSSOU8tLIxPaAG4UGYS9jaJqPnuvf1RW5k6G18MaWgiQS
OoCB29iztzL/Jr5j+8KY73tJTICRKq5zoENbYH359Kl2v8jBw54plLgAJ6cvEW+YIE5GY72DrxTh
Jr2kLLXihrvZMUE1CTuKdf57GvgaM+zgg976BD8JnwRkiHkRNNJczF58IYSSbOU9h9S7qYF6DIrz
gY2AqG8d6hSSQJYv7eZfXj7JrvpyKyTc24xfH9Xg2KPe9SvHiXsavwcD3en7GALRpUFUuRBDjJ0d
yI8TiVVmCANxrnfKePRBTBAdBv9pJ8/Kdv3rf5akKkTxRSgUzdjFZ3h1Invuj59yEUgolTss5Xt2
+SvWEyskpfHM808iHj3ErAD/lYoIzC7FKgvm9bTBffdr9YzQnhY5iWNBBLDMayAGSbTJ2OG3xM7N
zQqR1EuK1tRNMH/GW1q9TpafngSTWmf/X4hOeaw8hOg0XpZwvfBVWgE3ub5ow6cGmRLxkKfb/03s
t+bolUGZDwPcw7UcG8/K0nndVKFMnu8hjk4GC+PGe6dYmmgCOVTf+yse7HPb7XmbXViB3frKS1my
mvuI3S9kS/4lHGdMglADumCKSEALqQ8mpL5c5i7GfkTOwdJC5EL3EN3/PAHyH1SxXwLuUjdu3MMT
Gmlqk6knGAbHJ2mxW+d8iIVIqiEfXOmcPE5nxwWWG07k4KStM9QQTZr5Of8bjdNe6sGPv281Ix0V
2dzmKf4pf3/15izkTXbQtXFL4EkhiyMzC8Micf5vxeqFtEX+WC6Q99r3gyW22J1TcEvDUkMHzIax
9K5nN47PhX2baErRK9Ujch4vr0XlMM3ygPBAy8w08ZyX+/u9SU+nCwinSGHD+mr1rG1aTfR6TxB2
+73VwIlXJBAU/j3Awk1kxymWTb0EqpKcWbKgzrdyxrow1q/mmTcmD2wP09pC9FbektahY/7o0Jke
aDdS79Aaz2teBEKdUADDbdZtCkgrW7qPeyRgZ6OKz9bkRipjOPZqmyokPMXhMgdkKfdhneiTDu13
7aVZpTjJf7GKPcqUmdbOh11RuEoO9mWLI7qnZP4So7WNQNcB8zybufncxj0Cq2qGzREvr4oxCmrZ
Ivq4toumOQQowzXPGETWrTjc3zTFOxS6JZfcgvMaXB/Cr4jrjKKgxUmPOeQI+RQ+Vcx9NpV+2Dde
bxncur7R0tJ76vjtHuz7LM4VjNABHNdsdCkAM2rT1JTl6E7cflb12UZ01oTzhsqB5lmn6CC1a2Rl
U5nzJ9JSIRe19TfPGzaah2THDrBo+f3vAbfUiq3f0mDZk/osc2ZceNCptgamhDM1nQY1ggvROTa7
fwBw//bCyBuC9JZwO/spADqOhYTmNmi/z/E4MeSs9qz1bNL4BoJcbvLyHyXmJ4i66bLahr8+iGnX
euOHK3vmldAkBNv6B5BAZNRGi40zZdpII1BKUZ24VOE+ukVoBBl54bPbwBrRWZMBLxTcwVwM66zv
0OBzoDwTMxSoYMHEoIZXEYzGl0cqc3t+mA9vPw4tioiuV7Pt4CQ9jfHvCX/7SQ9a3xL2le27PxEw
1+zgjcbf505RxBL/dj+Wfuwa2Okjx1eM01O7l4JVVJVYQBNgiRIxHl0zXQ+Epumy/Uz5eer93CR5
hd5rn4ufYkw9hCzdt2a5ZtMq79/F2RaHxONkzPVhEZGa9BPBlVewJrXISUTD9p88XTPdPZaKfm5z
4vXPLP65RfWmfIx4t2c2HdwQLrc5M/ObfMVkhYrVJukBnztQ/quA67pqvhpgLOHJBNM5n+a7Xn3e
e9NIa0GzPYc0atkJRpqa9KYhGeTGPDStcVtAmEW/ol2iGLy3i9FKuw1gfbnqdoWDMZxx5PR4T/UE
jbzH7cDCgMAxfso5fjOBuncIT4C7b2A9rMgErhvLxhkAsHdNjf8M10a1nD56Biz/WhkUwmaAiQ0K
c7Oj8dDt4wA9CYzfqK/eFRWrNWFQoZuMJIBm6Np7LI+q4PJZx7ROuQF2UzX3r35D89vdGLTAbVHI
IBL07cBCCXAAB4Sl+WebaSzO8VG4eZA/SFdoaz9M4ANmKcLnASAF7PFulcNvwxWPQOBDD+fJCmWb
4Qc4n2OYqE9u4KP0I0CZ6lj4osKnshS3yLktXNrjinAU2v21UanIu28I1sPaIw2/qbUtypQsQJll
Z62JLHJIrAy8Q0mrwXj5OMWA6XmMs+ra0g0/X9gMnNZdBBN4eBvgwPiVzH8rkABijxpzTw1Q9wpt
7FNI9Q/LP/rjpsFyffkvut3GGoYJOiEiHtIpi2/+ccE+/A4L6v40Vlusi9ldjjU1L7ott8L3VOXr
oUvKlMkvQPy4kpiKCM4eK0ydqCGFM61lvLNhosZaSeJEn43VEtGFm3hHBRbutdii8iWddDQAUUX7
at7MMsP1DdYMPbP4gHlKlzgAsj/dcw7arLklFtkeDX9WlmcBMjhTCLp/7YNAr8kXZttTCv36csTB
xNdqE11gkhB45q3EinFrYtqj+2reiGR6MRAWuvalaSlJBqAq7U+jGB/+xf67AZalQ1q7aqBKFYvZ
X1Z1tGbOziIhRk9LMoY2XWOSrmXPBoLZb8d62ZTjpETp3ApwOSncZWgJH0g8YRFZU3daDohibnwX
lypeX71Vk9xKPCDQR/qCPHJG4R+eZB2pxYtJnZxaG1Xls5NfwXbPUHNxBxu8CTpz3fRuInyBzTkO
BI/sg8NJbLs29fRrsfUWwf5YKPDXbV/Ov8CCt3GGyYvppvgpOqMGPnJ7jac+kKiYUdcfSvTNnecx
wx53Hd59llHhFFRFAvW744gxl32pXTFtPmHu3nzgJ6+PQoPO0y0OGirs0rHWKguLVG/kpq62LfAf
lA65MFPLTrKf7fUIf+o/pnlQ0DWxJThVEBhoVj4oQ/yrNUAD2TJ8JVfTipJWQG6pdvjqfMmrFviX
FyR95Dwn5chEC/P+n47QsYcl12bYFWTF5k8PpaHXwTWGKoU8xQ6fxR4KLoz6V5klVEKBn0ob5JSR
sEkh9Cr4Zn+uBMPCl92JEBHd++HHZ4Wg8bKfKczPWmdE/mL9LXFO0Vc39LmKPJy8vHktQfuiTT3a
x0gX1MF0EfeRHKeOAc22BrpHTXUGasQQ4PcS+5kEVF6P4JhuJbKltr9ZyAvlILjSKsFpclxcGTvE
uDpo/x73XfVnr4h7yOb5si9vtO/+bqNuT1JXbaeBQl14/oIvHfPZ9wntbIOIZeFQmdFwAMtq0iT5
gHJy75bVOhY2No8trUwbwID79EMDnzWm3VwNC+oanb0uGXc0vtx0WUdSkFHr2SXORdJBTnZdiwG1
iIwh//k+STHp6Z0cklJOAjNbiQ0lYm7jM+fJ3PcsjS5vQLH3dB5TxdZ2ePGVs5eONeQXNgjlkTBP
wA7/qNfZncVKEKagbE3cj6lsKiKPmqPT/L8+5NfcQvxu2R6sxKf483tvtg8ikj4pu2u1yadcSYFv
sBzGLIC8eZe61N7iZgqk8nbwXmrx/o2UuqPZFbWM4TfZURX08dMggO0CkM+J7rKJHFzL6xuOIRQn
JbuHhGrsP9k7roNoxZLwSEJTWAow4RWjmYQruDIdB906hutwKnnluk8zMQnqKPvu0U3rKadvtwTG
KqZXt2dm/cdcq4ewJzGYg40DxBOqpXveB/RdI7WKeXB8HlN3y5R5DHV9vWqGCq50pC/wClqrdcv9
R0wcQ8IFw1Qxwo7/eGPiQLWIg0rhR7ROwER4+DzisgQJpwRTRUMtaSLdJYNsLscMs0xtTt4/aT5C
ovbNAMJVyNjeqxsfxEj2FwTxfoBS/9BTxamaB1MxSen2wwos9ksuWCSW0M7zTMHXlEqMvq9anGvz
Wu3FVl1Aqi2rV2cG/EQRdAgs3mNVAkiw4JwA5VYhmS7kfVkSExRiGHUiNX92aZGPbNPdzCuUAQ46
APKiy6r917nhYs9bp5zG9WZb2ZLJiwtZI4VspUPpCKD7FmHKVGOCh/bGdCkfAd4iTg9S8zN2Up+e
pinoSHpLDofkHaKJKvfzTgEy3R75Wpv/ErIvFB8xMhvyFtgIemMv3TehtFPf7xMh09OGf/ai/hBM
F0eIIx3uhTJye13XOnAY7C8bmNqQeYxwAHjPCZ7rBHu6VASlvnsj6dupqefYUs9/92sfP94nkUO2
zAsTpmT2kiWjWZUJAVDC0B33HmEsbGLUTyraDfn2epAcZO5pNhtBJUt7PmuHhPZhkOVjyZCpo2wh
qme2u1imKwDG9iWZ/vAlnZ7SVpPM+YkYxxq9/qzklSGbxgooWewI3jZrX68ifd3ok3o4GTZJ+ILX
H0vwhRPTZtagHYDRaTY27VcdrNYGGvD8ookwgMNo4UAAyEBKGOa/jOxmJhv83ckU5M+kcP2IoNDq
UtX9+Og5FBPW2rqBeGkPUvyKwFrWXv8sk78OBfMl3hpN7BSxy9nGlphnG2bbtfw36HIHz1JGVlNQ
FBy1ox7uV4o7u8eNhZHtP6tfVNeJeRRuK+craojdoSDUCGoZkwnawYxyX+wpt7uEKCGN8KoSektY
S2ckgcPVgIRf4gjkgaJzoSJoMgXVNqMg2Fzsi1kcENIZ6GhjS28smfSk7qwRVoNsYpEwnPWh+mJU
99tydaDjC8piHLSUoZ73OtBaLGnFfTfngBJ1qZj1In6alVk0N3Lh32eCGL6m+0Y4m89UGtNWesjB
K6gFbOWAFzPSruz6MOv8bbWAZDkkNlMtmFQRXjm0nZcdsgkjezTLAoKvluUwsmugf2nFAkOTeAQZ
PIMh9uyzMwWLrV9PPPT2fDuiSeBhY6jTOZCZYQYf6LMeyucfgw2UAFuCLRWnvs0J8oqbfFAj3XgL
JMoU67BPudcMJUIQytjcq+au40tLFtnuvfL1ig6C78P8MakYCx4dqJHHO2Bu9U6QIqFruQaDmzeu
BmmypSa7DtY4Z7/Wg+zbtdqS6tUnULfjLY7SdI4u+WnIgLFZnFM3qkXZ+c9iRXhLXFhCX4lzvenx
+sqcw5N3P3FxPQZ/XIeyZcv2Lhk76gVJJc47g0IIY0SxZSaGhlkR6WEhLIqvcO2+bl6x8ErxBeIE
l5hb8aK28xCOeAOvKv91/fZ09h4MHUw3yxE3IjZ4PLl81Yav/eNjuKH4vZ2NjnwaGLgnCpBXM7J6
wFmzQutdSM2unvlhKQ/JRyunJ/QwbLdVE4pRjIjKXN2Ox0KY6EXGUC8uaiX/XOTqmN8lgufR+olV
8zEG1fd+RMXPjpU4hQV7At7hVDKoejlSZ7pwQP1gqeor2Spt2jY2grNi9loZUA5zzyj1bux+vuLw
ehvy8R0HMgvgRwUF6jBpcB9T8zSkj3lEUnk7JfCSTV/uX1NJiU2NjCgg1n09BWTqcOLzttMletTc
bf3fdmGWd/QKzsG7oxaEc+FU/fhWCx0Ss94wXZhf6OGfbNUihcdQCx2sXK0pboyKyar0Pw6IVOA3
+aNxfxR/9zdCQu5IzHzX+SEJaUi0VQAhmin8R6BttHIu9AzeW8Q9tSTSCTvGCdFGPHf6+c2EjeMf
BeXGJnXwmhK0fM5126saYna+rXng+d8g0RywFtnmu/0+CHWkyq3JIH24JtxJ7sM932fDJfGFfHF5
W2FW3DQAfVnxdz70HU3BdmoxKiQTE4OrDCb4dfkGnGGhiSQ5zS7fm+iGiYMccWU6Z+9awn9racNy
NRdEZM2cWClHgJDEbB5qHCmJQDOmhgI6Q5jMUTGza/BJ9MWxzDFHe1C1DYBA+Gnqa1PZBkE1lQ8d
mO7/sVvXY4Ss6ZyGEZ4Ov6yANkcohq4IbKyCAOjMXIK+VdJplbHVy7yJlXWjlFRtUW+Eu6Z5YEYG
mnnwl00wT+PRbll3QraBfZ9GPoLNnWu7NHLEgddC7QR677T++5KmohewplZR2mp1wXld+Z9IsH2g
3zyDl2qyIuPT5Lmhf9pi8jgs2Puuu/Gu0oIuMQFfunQIgzstEDC5V+L0yM9+Z1FRES4i3MSiijL4
+anRX4JMb6ytoDi0rXmxeXiUG0Ji0PoVTcwmOJyM9QBmGo0bKAyKfYL+gX1KX8IcKQELR6nYKP+Z
5PO8APe7G6SOUYqn8/bZU4gfvOAbD3AmKLgdF9fuYhXv9N55xjMk7ly1tKryjqBO5rFS+56IbklV
CXmzj4VnLMW2/naUf28R63Ro74UDgQMy9C9kmXmXDQQkNlRw8IKLu/53Q6aRQWCKxOzzY7Q1ZrR7
CuK5um2BzNtZ73DCcWzciXxdv6pd260Ct8tqNkGJ7Y3oKlQuuzkFkDb55JXfM7oBpqwHdZhu42zr
qePUyuXCiPAyhteXGqpoKNuv0tv6TIxUvx8GGvi0SMty0PoEha6ntis4ZqXRIe+qF2R5j6pGv2lb
wl5opeW4DBk1r6S18mQQXSva2l4XaL+LZf2S7AiBZOMCw4v1LT9SRqUPRqGCGCYqDy0BQx3BKYxu
xxChv+adJdcPNo6HjmCTAA4g/TmsNK+VjoZXmJ/6k0vYK0TEOGJ1Sk0H+4XFJIIcnJzlw7X6sJYH
xONZyOh87eMR8QnVgjPfxbQfMOM8ivCa7nU8kq5j+Y4oGum/V9X93NdCl7iglLj86XaTJj77/t/E
Y6zpfz7vJJ6gfjumBELNZBNeFCT4s2rm7Eqb3nZXS4ErqFsbrKnSd+bD14cqs/JYk5RF41g3R8gb
oDXEwOaVNr6gBfm2PRvrC4Ph2/jiGROLZYZmgWodwK+3Kz+5KdTW8S83T36evalLuLXijYwJDrE+
g1kTlhVpJZK+TLFx+0+0nMFNJL2j9H4W8W2fmB+NU9roSiE3j0NXRGz5d+motBrHJgrcAtCwkHIY
HpSRJPTEqcD8XPbPpTvO88ybP8VHKShd3a1RyWND1it/98I+II6mvDcngwS8aWe22zIkZ0Hejy8L
YKkhFM714IfAcVIlrcF/KK5B1QsxfRLV96f2WjwETM2W7qGM05jTRkyvB0tnXqtvDMOw06dM8GA/
A6C6m09XEA4srv6yjAQF/17H/vdJoALxeEqhh1WeePu0UAR5EDwI5YPqHoxSgit0ym913ED/7Wzr
8grBXUu2y/5s347saIUmy4sWEp3/hW8CaQ19ec8GH5fLA++bhDcM7B87eNpJl6OlQU3dFPGNEE7c
xuAt308ShcL3HjMsEJIdhzwm3UB2LrDRQfWOMSSZ6HL++joWp6Yo3I5Ejt+Di32bftICbPOaVm2n
sb9JAlUO8FmrXGDdaSjeiR5fddwEMFVhvjOPcHRElikh5KjRbTV1e8PV0c+A+jbo1OBK1JlFihU5
aZpQokMWU+KFLK/TwgNzQwAa03pmN2LhAXQF5jLYzzQsxuShFdW+zqri5t19WL7ZQCojmzjokufU
ski0i0wpUa9bc7TsAPGHYRSRmq855UtundKVyenUAj3/anfmutpVAgnI13B6H2Un7Kj2yJUsFz/b
GEWDxK7xWP+0RQ8YIz9yQfDDN5MLNVCPas5xFl+HUDjFnEO4tGH39zdfiQDlX/RwCzxPrfzbqIyc
o1YX4J924TU5Relwcnh7MsYEn0a06ovkhRklMYn0JUD2W343Gz/GP1KyGTc4de5AsTH5gHDPDwKE
XGC8qts9UzkePe2Osb65DDCSZ9Ort1AjNBoHYGxBCeXq7NWhpt6LKbVTMws2VAW2dtF+/dAPQ0ON
j14hDm04CZwrF4sf1fT0fQMDyAgfdmjhkAcozkHN+w4MkRKs6keN5SCvp09G03orySEFKCCn1pfW
Imh8MO9hFcw09nsx3ah6JfJ1ofoQhpfUSi/Ea/pCYQFWyW0JyCTfDYVLGk1/JimjHTdENnIo0yLk
M+BnoL4IoQ+b5saaFHQKzWPqky78DpylIaoZhdEdmh4ueXnqMq1bBkw65N3eFrmviLCovsLrKjvA
Lm8xFn9sCILJFUsck4yIuH/ydEhR1TWPtsekNKYzBbJy544NOHB80LoR5luDe0+9cVnThhgVMIUd
40Tkro+yTEk+M5sq+R+6sXgWcosXdGlGLx6aTjDntwGzkBYR/bVLdVwpB3jSTz5CBTHJ7UDecE8y
RIKXPQZpSr7XCkflMMu0cxUvFlOHcPL2z/TqONwTJ/io73U1LXyhmnn0DTYrIjiFByJ/kZ+ZjwzG
4sV1W4VyZOSpss7KxWaSqsHh0193oFUgNJJT7M5mckcZ5yVPBEf3N20jcEUbNmPQuLktXwBtpboC
SRNRmdge0k5m5/ehXzUS+NDomynkNmZwgQlcAL9l5r5mnPDHVuzZV7VfFDdutq33ClFuv0KUIPst
keNXXsp7CkH3SUZrmN+dZMMHKwdcz2PsEgWNVFLz6eOhclgD6yXoDOcgWLpYC7UrMW+JbaLMUvnn
N1pv2OYtfyeKDjVwDAAXdo6dXKzGL+befUaF6Iv3/GVmk60V9+wndaE/JafSFPOYAbmEh1Y6QcdU
nnBuOeLTEdC2XRUJssAACbP+6e3wrOclpCBxny82nw2Fii5A6l1+kB3B1FsWiNL43/TYjnMrwI6o
GKxl79JOvgycuOeA+3LaWKP5ciGsztViX+NKaMmzdYFMeA/0ECaLU9F246AIVfoCGxx4x5spkWR1
19vi7IHAKYPqbr40y2OoDw+c7SViWhTOusyy8cFWfSsFvlnz90pAmPhTEEG9e0D59F/LM0FHJWsj
yR8Iqzo1wsQ4Xj9Q2FfjdYanWLw0Ff5HpcxzsLN4KW4h/2WRgRnQu1muW9+9Xkpqr3G/zysYfASW
FWGCgw5tdQUhL28KGptTc7NpOhTYB3o84yXJ4XKJ7LiGyB4SLRxUnkEFChH5PQFDOUHUINDPPzBm
2JOG9vIVC8yPjD/7exVkf71qDvFyd68a1suPK4WpvQo95LuWWE1ckIf7zzFbb0rBPO6yPNoIzOe4
XIkV0pr5V5igGGubvyBAYm0xKJhnPGHSpc4diXrUzhLYP0vuQp+ct9NWspJUtZ3YvGw0uArClO35
O9k2snHy9xD1i0FoYCcBdleLhVB1H3dfZNiCzuJI9fjXo3cWXvvmdj4xwIgbI+rOrdqdo+5AtnqF
7sTyIdr9VQ/Thsc9sr4FBl5eicR6Vgfxg+pWiGlTLfmL0aE7rv+s7WfsG2sSLU9mJOGQ6ns/1yLE
tc6Qz/Qgxv32lg0HLjluIjLOIvF3HpdUPKGJ9Ji6IUuEYd5it4VzPzE5AM7wS4jSc0/SBNA7olnE
6fhYrxKR9fNdBOkEw+hlCOSiN4IO2w3en+JWVs/VUtQkI0UMA93LuInNhm3uiuCAUr0Gs9/c8YNV
D1CuQoUzH93xrGo4BADI7j+YF1D7AN6WJb4TDessJ5bE0qEblYiRKfKxuiwSqXuRRKs+qOWrS7l/
s+T7THWjW/gsu0AJb8C8tJuuiPVC5OkIJ+xNpnP3ubNvJuoklFkCgjXvKNX0gsVm2Dke2CT5KDrP
K5ttZ75HJdwB19H+RMnf7mnkUiIPIkUk/O4/tA16fGUyie9zp5uzUFxIO6Ynl6ad34O7GRjxVkWC
teYH19y3Ilf9AKAiwhZuABdlnuA4yyTo9igSWpf/LzjvzHwD2cafTMOxTzza1ZOE9VYDSWwGhgft
IOk0iBWSEVoV7ZSXsQB5u6dJyK+Gvj5GyShszW/tyNyUua2dBu+mWScNqh5icY99uAj7N6O40uhZ
hLC+pewhXZ61yZDaOwHyeRxYg1yDAfYT5KRBeWfiNvyEeE9lmGmhpWl7h8YwUmSzp2kb7kh+bNFo
gyVx63ZWTsElg4QAplCMcmmx/55MSzIOqUJNG4BQIllwJx2OoxslHalb8UlzQNjbvJjLWapGVjWs
I7zDHLhlBB9TPGm5l0yrKvYP22VMNQjaKI5mxNlqiVaJ64K0tlc2lCf5xed0AOnZE413VT/Le2K6
fS8KCrE9FlzOvkyzK+5ulPn5+74ykLv83nOppgvNU4zV/VpvzLnaqMxlLu21DLk6tvCauA+/7eH5
+uvtEOyaLUX1WE82CK58dnAswrc0e8/7oa6r8H6g6fUGoG3MumOPVa3PCJuAvfweSKht7dWyHJd+
nm7VzoAHQSl6RyiczS1Kq4TzPwZ1aNDdOrdMpCFFshdeHvx5lfhAFgvfJ6wSGFy0AzLdW52gCsoJ
das9hmxyOnqk0qC/uyUi4lbCDgSSdYF/cWIkDHv4ssaT7aPmUQphqCBrGiMeuETblitK4L4fzUow
2RH0oUVOj7F/yj3kKFrq5NrmpKPRdW1sdeOEkKZ/AvnFKqVY7yM2kNY+wvqFkuGbbNK5zrRUgGTv
k6E85kRULwaoh7IDJWyhY5zeZzYpt9KFI/blrt8ZGJzFpwQp5FJDpHkkPLJIgYkMsJUeVMPLWsf2
IX4ZUmhwlfQrpB+yxTPlJe0DUUDTW+sC6AcOn4iOa/DfgMbOlRzBs4kfsgn8xiUB0klBJTicwhIY
1qk5h1uxgaTD6HV26jqXyVH9pgBbvKMZv0iGwQjsF389CMULEf9hVpE8zR35Ah+Q64VM1Iyhbea1
v1ikb83RLt5/AY5yjVyfo0yrvOXzjQvaakucdk85fQwulOKVqbICVjRJDVoAj6QwQR18gQl84Or7
vGF7GfFV6kLTN0c0knrf4xsWH3i6qqAyRaCTwHh4W1YoDohNUrg3JVOa1/QsDd7CIO1wBpA4k/JO
Q69t0jM1lpKCbxZX2XcMCZje9y3Tdx3OwBtfrnrIIhSCq1abgfTIngt2BjGyZjnzYFvJ5+Us6WkF
ZTZVwwl4/5B/VZ9DxEnabD4QpyJmHKODuJcMzyoIue6hPTox5sBKBZKP5gdT9XouyuQebbGJ0cQK
nvit4NNITpJ4ekyWBE58k/Dl7BpgWQArraSqDYlKrZtmC9832Tsy7VhZyi/fTaU93HrYtg0hC0BE
4UBNND4GjyjuqJKg9nEG/hhsuY3Ph1F1gQE5pm1+3HnGMydvrrVA4YdDAr0AQF92bDGSaqu8K2Bw
7NB6ZMm7Pc1REQolSg==
`protect end_protected
