-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NlyvL0CoXBRbsOmRlDihIEU5UHC1alBGxlHKc12Vf6sGpiyc6BDSW61+9GC7zCMCHZZe0tqfNefr
rbZWaYJ+D6glkFFdWodGe/FLPuShRjrIbEllERHv1Pq4v7MjXI+CyLj+bROXVPVJylR8fJ0CjD3N
TS9ibbjSJgqATi2KICoHScoj86W87BJZQOIWNBGrdGGtwemIz0G0jLqefECG/0PETXuw8KbXeqox
F7taNaidhStbehydmtgGQki6tiLiMiM38HfxdkqM2pWqID3qP41UI2L7HXByeIOmb2Zz0I6P+P7B
+o5fPJACjVoG1gI9y98PR/7I80oG+9bYjF0kpQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 83312)
`protect data_block
nOXGhEkI3QFCXJNn29Vj33JuD5WGolauOEvcB6ZYwGUAHeFwItTmLvXN76flWA4wVNMz+si7/hbM
r6jgO4eSS9AGEgQvpTHrDRykG4yage4jIoWT5xAUfC6TnFjtly4JqgQ9cV0+BlH7hUjLz124+EJ2
/FJ5PGrcXiu6+ZM5r2Nk2YsnQIqt/qu6aALOY0vuSf8Z3AlnOH4rJZZpVb0hgdLhafh7VdJBt7W0
Qcbr9U+FkgjocLV0+nUtz7xIIeAoXT1upql8gy70zYZzZ5JdBGe7aw9FglqfwccbBZBXtr4jb4qW
vqA1a2WQEiYEn4aGrJs8Hec/KKa78Q69nYkWdHDuSjLAO5NX1cd2rAOBqha+79FyvldEOmccFx8a
2OGjr+1puyVe+n/WMsowUSBn06yMmPgilQIiTAEDABp43nTpPRWJXyKE9iy13xk/jQu/HOx6+7l1
UO7GtyU5ehMTV0xuFce4z6aoJ4hWspT70d7frmNKTi6KB7OtE7y1O2Kerdsr4ziTDIU1WBD0Lr3k
IhHK54mqCImtoFDpvDtDztX+keqXLdRplAr8g8KD6o6dO8kYELdjVXImRe7459kmcA1fh61nxPSw
7Prp281l2Lc7m4HX0D8fgy0jmfdgw0F6qhK4Nr4jryKkF+jyq4hzm2B4lrEUZVQm8eHDPfoWWyPU
BzSwPR+G9KfACePlX5KiwmWf8Cr5cf+rGgIS+0TXnBsjGoBgFOcejPnZSI+bppNE0DBevyGM5JCt
TcupA1tAkARqregSTsaoGV1kXOI7eO+Ss4FAldCw0QJ3aXSUaCYafdrroIMc6uicDnrN7geQTjGZ
i2XebZlbxgOIAoWA3t1du6WhaoKvXfqrRIz4gt+cKVmuDBUyunkhdaCB7qCW+m9CZg7FWW4pRmDS
6EaqgfHdQ/qI++5hTPOiCxt6n+nSfA7/cQqlIrWokRzyp3TVT0ETJWv6eDJTHt6gsbfbsYEzq4ZP
bYFOKZwjMBgJKQF6p2jj4h117r91BETDd1aDJp/etY6u7HTxooo9PGjiVWRF76qJZlWF7hS2KBAQ
qputbqPGK52AbuwJwy2SncEIFD/wuGX5Wqqx920RUJIyIdd4Us7IhubEVKbSpvlia6sVv6IklH2k
vXWQOauIOFA7YxAopDYN2h/vit9AgxTJiyGBiSyacyy+i+bBeuui3DUsm4c7jkW6vonywpz8M7G3
USWQcmkfQ6vlyjVY1MzKgbC5l63oTcjOYqSOTjTHaWdRc8Aw5H0fAQ+APul6WKqJn5EkdkVN/sJq
tZ4lA9DFs6XVyAf/PqGVpy4iN1XGVqffNJhWrp1OKwmKILsxeIPprFv91YnlwxVSFNqBLyMxKOpM
NUa8jlt6x1vAw9RJI0k8VirklchwdEy4OHg7aAAYyfNcAJi+kMHVnNT9vaBYiNMjSWfQlRckWvVb
mosQQJZvGE6QQYzd21lv31LTdq+EI1pMRP0E5xoUwkTP51cs4JLJMVnI9Jmms4V0SrIUSZgYgrVt
d0+necYUtFzKHov+GmGaeN9qwjOkTmjRN7KLV7hIuN5RBN4eclZGCIWPPvfQwXzG3XS+3MfPyKwB
buGW8K7YD/t0z24pS9ZRw9HhI7e7jU9ONsM66phfpFwt9l3lQAZAi7kPYIcjTcCR2Ee29WhjKLRc
5CPxrltfPLeOT//RZx/oKMIHJfxN4cTzh61H4mRMPU6JU8UeXYBQ8SIoUaFLMUGRZgE2muTtY7dH
In/TLqYxM0VMDCxNQIxeIkTgRPvEBxOjUcG91TL8ybeBg/l+wRaZ0UAK9nJatSTFythUym+skqUt
cOpwjDtg1esQPsHix8p+yP02V4iMcCTuA2JjXiWdziBAM9RTt46xq66ABJIIftfspyIKPy8XRf5I
TQIZmKGNASDK4Roigwl2uAun2YFU8yWdJtqWdZYuG7y5l8+F+LF3FPKj9LD2YclCJRcVIpQ3F1wc
xQpdlZbhS2AcEtK2aw4kDJ7UnokyX+yWz1U7tKBjILtO/XvlDwvL5mn94TjAD9TMYsMBnLd7bU0s
dmn58huJMKqVyZC0kNH0lYULLqPVSvuYzJ7mixyi4DgIRwJTeYtvdC7QVWIuk06MEHzqQrXH4RYB
UhaBtxpWyfKtquPdv3aSUEtnrZk3WjIJgnDrs81hnftQtUMs7qlk0/cA9E+Y/D3WO63EJdZx8u29
XpPc2n1x3AtHZ03WhDEfFYHdvHXl/fMRqU3oc7tYl974E619ES/pDqFnvJoLfWoC8GJS5D6JZ3NX
rlWZzTtFkupgrzGxciutQBQN8dRNPkuArSoeAw17ST+fiyUfT5vtynQt7FCAHVn+2qmz7SxtndnO
f9XePkYWEwB08UDWbkFsueIraNnmv+QN9HPH9QrlJM7hK7OSbFQbU5qOphOp8RlzQjnPF0WeI+gk
Epp9FFRODmAEjYwPpLloKXdPYsYag6+2LHi49KGYeV75xaihUzvw70K6+2sUFUiVU2pKWpnIB1y8
1IfkDUwPPZEAMh3+i2rYET1zF9yG91ktgGOMeI2tDXkU7NitmlrFn6E/nJeLY5dt1HeAcHcYQ+FK
/PW2OwLMr7yh8JKZCjoOZQHKFerlVslrzyaiYUb6z+OlDmMEVw+Ln8LHGbPb2OVbYE6E7iYWClni
cQVGjeGwgSxPAWdG62ZQ9emS73+Kv0ElGgtbb/lq+dJyeYTbN1ne01bLcG/fOCOBth4ajvepbxPl
WTw2Epg6YKcvLHAv0LspUeUYJuzGvkWd8nW+Zjvf9+XW4lqPpfHlsU4Wcy3R5iK5mO6MCMnNfBBM
5UkFf7fSkmQmoE++SUj5+n0XdE64M0G0KPIOhZAtnCPan6abeIMVlPhXVRd74QQ7kH7ViIFpw8bW
76a7MF4OUyQmw6x7GgspqZezwQm985NBFI9bEBa2lUJVa7GgAldmOfSXC4UrRL9IzrZ9PToMTDuf
1fGg9s1VEs+R2bQflmQSD8Tj+1m5uxdQc+A42gl+/szCEZuQbjNIg1Eb/kmCBPmP7mgpx84y66mY
OK3Y5/mMYugdE+pHLlzpLRFWMhHTBgenaA617PlHy8aRU0EwxhCblWwez/o2vb32xg1QaGJxhDg+
iP26yoCEywLhRDyqG3Kx3LF08kQHCsugAAYJSvxeznw0xBjY8KrvNEt+WPIW8Hbw9jSpJWIzO67y
UtwM8YHo9QGYqYBQsIivMxpVnDHSigeJ/k9xSD1gxQ5HwStxxOaHUDtJr1ETb/4j5teohyw7QKPP
qSghf9M4A7q4Ie8qJBBb6gGXgPnMjOf1vwqlhf2tUPmCINp9YWSfCfTIVkc/c4L8/6AIOF3BOKJH
jpMD07br1Hy7ndHJSjWsYm5NQogEMSCW8dKDj0t9aGMg/pmY0ru0fllzojrJYfMkTdIoE9RnLy17
7FjcqudQlyi6pEdJI9afZHxf19j3Eto4aUZfURgtza2oJ1mJ1rqL1mlag0MBDIVHGs2TbJ2+yWlL
vqvAj/O/0bp03xt1Au5R53OCMpxSrxzsBvKoXLtbMg/Pj/3SM4n9htZW+QgBxsbKaAODjkvkQXUm
CwvL6IbQMR6COsJ2C0eTlFWYUFUvHgXsUIUt7VC0mFdKUkVdvgqfEgvwdMSedPGeqn+w4LPRidD3
r9APQM/FTamTBv4/DgHiXpGdoSqOQRNnvDIMh4dkdu+cmX8ACGzdeMu7CJ2DavPC43nldtp/1eMg
barLvkxgzisvcHWukE0107ADp5uxnqhCq7UYipkJOM9dEKSe6ZJwYo/kVrel0vAba2kmN2/tqDGf
CFB7hTiP658Rz3f3kqrFVkRLYuo+tKi5wzY3IO15PI0MKFPvyHL/S0g/PRdwOOs+k4+1N3wV13If
sj5oCWgs1RBSYxxoPdiIy5nPS5lSaH74E+3EF4LF0yexA8Lh7nfWcaiW49H8rkGf5xO7E484PhIQ
ZwKRWWw668wh1qWXD1Cgn6a5EZ2Dn8vUm2ecW5Ine3P53Rk2zjtdsOisvXsLrmReldFm1u9ixTUv
VCCnD4nGbMeueBIdpO5IxK62H9l6wrm3ZWvfSuBU7clic76v2lwJBaPgO0oFvxuRjLpzb+joD46r
8+GIyWdayjpjy+lXtUe+7nkacDYs4U+w5+JYdo5dsUDNDclQsm1+LSFac5GfEpspueugxlmO16Gz
mBxhUEtGDRdEfsTcqjHvZZdpm3ka2FFZfuPhUSNiRhKd4RhIv6Jx+G4DTpKZo2Q/NXcuoDMgIvch
yAl6wKxw1Txkhxh3eypyUXGcNqXWpDXBnMzq5lXWjdnpEX4TAsXOGJ/1GZpLpxl2T52Gqv3WiZ8L
1y9wsqzbaMy3YLoM/O1xuLsaB4BE62obmmFP+NHaWTO9WQeLr1lt3H5g9LyWvMoqXA6hnDh/OHb3
BXzNtnH3enkqta5U32bFbIjHlNsOIgFXN5Dxdu+6UcMwpGLoIpuLgoVh6AAeTl2qFC+w7gFFSHGo
0j7pW45w3akJRyFUqEaGNMBc+1EI5gH37bW1qQfI1jG6Ei/2VoKvUXvlnZY8ar8cWvQlarXuDxBa
FFMnC/ylTLJXarVIAOUYC/UY46S0aWJL6eS+wKLJb/eKn2El2fdgGbswmzPCZhh4khi9a7ct1x/z
ruumxfZ5FT/GsqsGOcbDqGf3Qn5WfRBCIk6SsC9G/reqXIAB4gnh+HuPGzF0V5rUGCrsUDvoRYXa
Shc+bzAFWI/7Hh/aF/j9KZa6D4yE2Ek9DXfjW6N+nUPfedpJLYpA/CCuUWDWT8co9ULQOrZflntq
2ORAooOMhg3FPlBaamAMzXPT97bKvzkRPAHSijlzamMgaiTs8jMxtVoHlo004y3KpTdMNI7ZCnEB
3ncksf0fNHn/e5c8HWRunSR0qDb/JKMqT7xD47ThpCag9KTySebbV659yXhjLvoaWwf7PNFnkupH
qMb2kipyfQ4ZmVyGvNWzQUtPmJdrxEoLNHNbg4nqIW3cAiUy9/3yaMLh2+P7MDy9AAUhdj92qkRL
6jmz+CQOR1uo9BOMLT5Di1/kgWdVTGNV8wqxPXAn2hJB1J9YsUZFmLhG8ff3mLjYdAb25DcwngeI
xlY2d0nLfYsfBaa+pKEcCqkLuuZgcwwcbyT/7j5EtCVqHdIC4O/E6WLjlINIWms/IaNSEc6Qo4s6
r0KqmHkXPt17GQb0EI/QY6aSSWuqWmUsqc7oJgu3pEk+XiyTqRneOnMOB3pv3pHAmXJkQl+AKo6G
OweS+rYvqjd7I7im0BNGdcXKnL5osW0/9xmvqoNatFaYDHa3PuGYrVxgXMXjurRUvRbnCopz+Gkf
GrkkAcWOv0p5zy3ersVLXivcwhScZOH+hIht0DcRtPMYBV6SXdC4Jvb2eKDeUIKsPOdubD24HQYf
7o/Wd1CdFK/mPWd2hOhR8Dj1JpjzYL5Wwf+ZzXjav6oj91MhhE7rqBnyTIYJubKdosuy7dQwMeQZ
k4SshQnt2Dkf7xcw+kdH9rAMjh78uhZ7p5GVEW95o/NejHoCJpnHbDro9la+BkG5YqGcFaLX8OLh
6Z06KEeJijjmCPdAgxAeYkp6EbD60R+1CrNs6HH8YhBI4TjZ5BG58jrpqbLjbRgYbEk6Oy5npvkQ
Fp8KuLch6vF40N7HAP1K018JsvyYhiNPElQk6ngbrzZfFMplFtPbf0oUDChcvrftQSPHH1dec9ax
rmxTbnhJpVPEJAz2XC9n2ZeSi9JY/t6T0TWx9ib7kOoMhL6MZ2Jz/3rydPij2gns5kKm8jokyj4G
b6EMInzIWpmnLtgj09iXk5S0JvcyOw5k1xD7vyj8zgIvDPrGNHRkFGg8b+qcNKwA7AkXnw8c8U4a
xpH7QXiisbLqvwTStrYWR++JInZ8O8VsSDW/3PUN/1UsMb4m6KwrUgY06W0HhY/FHa1bgnCdl1A6
L1UT6oVGdH8NmqFVLiVbtnFj+dmyyWddIy1Oup1vvg3WRD5An+Cw4uGSwCsA5ISR1qkNjBIG5vpx
0F92Zelx6BsGZpxH6k7RQVkF7/q7LoaSoBLKokdkBpAQiriASuAeO/xDYMks/KUzTzeBGsYMyZyh
lsvcSa1gzkdAR+SdHy54IwH9Yo7k6hBDLxgVo1IFsyBAfdKLgczdRdaJWY/F8NDqu8rqXZBGeIjd
luws1VGcjO2j1or9VMqypZMQiGxad3mdhl1Sh0WbOcyQjUtyKAZsTPOmodeRkCrphCEiTRwL+fX7
YstizBKMR7tT/Jo0arnayc9HVy7KBut4PI60Il7AHiiTVSYw+uAPHPCvlI5BGSIIKnweZ6x4hTKD
RX/umgU9V5qqOzNkQV0FulmU1C4VkXhHwTqBI3Js04zZ4G+QiGcboe599V6yPaZVhnR366NYbZ4r
jfOqM0clENk48iTjQWZqhKz+Q3x3PzJyKI8pq9tRn+Hr1000seCi4gfe+HY248G1/fhrFXzK6Buj
ingCs3JR0Ee/oJTQWjYaLc4bwvGKZfWAgXKbyOePl67C74jnVBNC6lI9XLPoP6pUGl8UvyhlLQY9
n2neMKSlcS080KBBjT4WHfLQfkMlHj7inbhXAAFiDVzrtHXSa+ByrlfVtM5r+C/feGzllro6PpJK
mPaWbVYE89uEqWTTYEYsg8kZNpOTxUbCDH6qjH1UMjV71TBO+SqQfmbTT7l0l+gGfwbC1tqluUqQ
SPCxS//b7/ywWSAY+HYm3DvjWNvyqs5PwBU1wnLVnVv6u64Eey7wPB+DY9yGBd+3Zlgu+C0/u6tn
bn3d1/Pb7+hZ8RnYoWQhNzPzgEbAGibcyzbAPe+T4vNcQD2Sxy/1nN9b/JdYXXmfMf5ESPDpkRhK
3NyYCHvZWkURzWmURHC4DCXVMvWcZYhr5NFBzQKyfv02We0zfusGfLB9h2vUwh842rqyp+OGTvBc
3doo1BGq3Wfq4UkkYyErk2cGJK4bcjKdlEkfh3t1NsLERQHWTCgvinCbITi4pV7jC1U9PBa+3Tx5
Oj63/W8DjzOnJMAaJtmWoPPiruA6fk3Yn55rWJJ97EKplF/8lyEUoXjuEjfyOqE1+gvBby2yqYXC
LyDMiWIALSbXLcz44Af41+tSUqtwsRbXXFaUQSm43rrsnk2Y3RmKw16c3RlaCQgnxNxBS7AMHpPI
QxiduX/YukqDZb6+aFs4HDpwuOq8sLZJlfWHj1YysaVR362omo7SVMeqajGdHp9copJ7LM9fl63V
WyLTzNGzD83AODE8J9DZzGQLryv7VXJ5h1wDockZMhYcr5vLgi/+/+UQ/uFZTB9pA8NawQuMOeJt
HWvg7+ri9J+eMEdilteKYyESw7PtLcUb6AbEzCtPANO/9esuvL1iTqQrJzBhyYID8WAVeoohZQ3H
KPGh/mzEeg+fNmEFWpSKmaLAsuo/yrOCmd9jOxzigYE/Ft8SRSh4wwxd4DeKFHote17xM4wQCE/H
fZvWlRPn1UEVGX5mXjaXIqdShmcKOTVNS5IMhOo7RFvcQtGhH7kgQZmbhBLYfnzTVSZ/sAzqlcjq
O7HetziKe6lsVM0hLlY/Q/4VxNliUdTy0gu5J19dfPw5fEDzogn9YcuYWV71mnBSBKVGH8e6M6kU
i2IPqxuqYHMonzFa1kQ0+fs0e0fUDGUB5ZS/aZDhmKrux0L2vYP18sACbuDhTIuDsxKrnSKXX0jo
2XFpGw28w1M9JR6p8oKHpvPbc18MJzPFZfNzrMGUuREnsnJb7ZhPGV2Th6enXx8fVW+HulYq7E5Z
S6OQMnUbB6kkEt9ow5Ze/WWmeaMhlDEIBZm+GMqM8TBQg5TR9cvPCVrrfXayfh9QACtRm27CTsrd
PVEiDswEwowC9TceuvantrQ3fVzAcufIKapdIukfJS8KKyIfhtrabgFsxZ42NDFMzp7yO/6olf/z
SYcWgJKSBCjB9VcUriqzzn+0lW6zWB20xR6FD619wBf/6ywImzKOkcmvk+Vy7YHMcLjrOjUNmyGl
XmxBIEbGoSP8IFZaKDzBZIzUG0JmPxe5xPJg5fUBsssLi3wk//a1D9Yr1QEgmG+kpSdkcY738dEy
XnsQ5+bQW8F6pSPjlvnVABXJCFewqlIBANU/bVsdAhlaE+YYAksPcfUrd7ITsxLNtEQV4lE2NFte
IX+nj0y+PocEEDqyfzAp0VReYxBWh+jlFIDLYduXqW3LwV4o3sl/jlmly2wGzQxQu210bInVBs++
zZmTUjf0I8aQwXn8PqKU+QfcqpNsWqrQLeTt0OYu8dWr3ewai0p/2bapmvfGPyy2SDpQsfaXJ/ZG
s6A6wqs8EaVrLMjNjDY59EKuxZ4bF1x3P85V7yPckX6SJ5628dYR1zROwsQKYRKONFPkSMpl0/rB
tkIH8GVXU4W8DIhJSEVtYhS0wsdbLqVbE2XwpAEbzc6+GGP67BrJPbVWuk0AZQh0rWbCR9G5tmBy
eonfu6ddCc9Rc78wkQy/Jb/LB6U4MDX2rPDjFuuUwLZBxj3jGxvRNpBKOs9Wn/VaCl5MZnmgq6EV
Kc12QnODgKu8o56gX5PXlao+fYzgwdeH540GImh1d7tu3l/yyyi3/nwo2gtsXOYwDQL0EetGb+jR
V71KSIEaiDnEVAux54ZNqTlR268GaneS/rMhzSutWKL1H+DqjAAGH1Ta72POFj26vEPu54kDS8KG
Z78NmgbSgeaMbJaaNycYalkh7pyYMppqYAh93EaTQSF1IdwG0ffYUZTFwwzOl2fLjkXrJGAkfEzH
1hQeSGu4GBv2oGTJk38O2YPJ4C/tSuV1JnihaYO95tRtUTm5uHpqPuZ6Lr07DS1ME6F75dJWVuwz
ddAHDhjq3mtR6/FEJMCG/+bOgnpDLMMOPw6xi72SA1rkrEyqPismNX0MNIx65K1xhfBLLKG6+94s
svUwHg/n/atDsNXCxYh3b6t2mkECzD5OAAERkLQPAHjIpxtcJtIkkIH+RwD20DjHGe1nykqM2+HK
chkcSoCp1+2VAoyFLJHoULUfB/VnYqL7xlXt0g2ALREIyb1zUq5MTLPgeYjF0x4eRSjD6m5yPu1X
P9U+XiQXTCpLAh5FN97z+5haykPKw9T/KFELOLWDUpov6cJO0mke1p+jB9loUZtI4KhU0g+Cc8Pz
iElpg4LEJXdaovg9mFsIEaQlsObPtSSfGkaNdL4ela+RVkyk/N15J+RVJ3pu6ptlnC7I6tcTB0Md
AnabZyHYMdSTcLGVJu8H6+99Q2SJecHHDXb0q3sqJCelcOaGECWHrGtwuVdCAf/7loUdl/nPlF0h
a3Tg0bNSsUgHVCNIGEJxj48g7iRokA0i8NTgjnwvuG9lekTPLK11zvrl06bqn/FtrNnq1jf5O74O
Pr7zEN8cYbMtdwb7l99q8bT/6A/nfgtutTtZGmdARRg7IWuXJ09lRcM5mXnXGZ+o9mbqcReJw9ox
A9nUKO1w7ctJxye7oDIRVEeI64O6Adnar8vSG5KUh8bEc6Nal8bCxEp50+5OA90G6KE4VdQnQQhd
THyQFWKtNR7RLDwgLL4o1hNAhtyXqZYBvU58KSzvRREYXZdseb/BizBQfSpvuKGLgBLZSgYPBOXf
A5uAqXPPGQrzpydkBZA/LpUHoiAlL8EdM7lHxmETVTCyKn15crHOh9K5JzBbk1gbInZh0CB5trs7
P/NtkvgiLDmXkSdRKnxJWyA84XK/J7gXUO9vo9G7AYxZCT7STV22NuiYRitPbo/l5UJktcVv6P8w
fdZ6NSFoA0btacCet5mpe7RrUTo5JOPbnzbhzzvgjCTE4uf2F7HDMzGJQjiMIbIV0Af99c9Cl9aa
6h6Nvy1CIAZ8+Hcqf+lr6TIBpEqtxZv3uRACHvxMmqjGp2KgNEl8owbKDmE3Q8DF1LSuiXQk31CL
lk9vIPGBIgV+lbXAid83YebJlmrnEtvDq2rbYhXwdcW0l4ea6rgjdxOVCYwPRm0McN03KTJYvarr
ANhU27cXLJVCVSCZjmIMTwXzKNyglrGaeq9kkpIZrgRJ/0RJZapnQXXu3dt1q+GlyOltVdt1x9hl
G4teEBC+u/C8XmLdoXdZpynBSwKH+cdh3vgPRvr1YzQW+hSZg9UhO3p7Xbea4r6+73yzls6YUqAx
Vdex3OcNID3D51nyr9uddPxxsBlpSg0+kjf99ahEKj1UNZ3bny3H3ys2Y5TB2YtqS3+RLNZTFGBY
4P/D07tSagLb2lX0dllfNn/27dqbMOfNA1Hx2Wko6qOvV9yvxxHpsZo9wlaCkoxoF0sxIKOgip/X
lgC4u8pa6Pd7XFmkBdcNNhudP/NUpqXAnhhDkQ+Bk/p3vJtjpMW1gsANt2z4pL4XaZeP+4G2F09c
Fgpz8C5wHIYGwYDj87JDuBwGHW2TmOALi/rIyi5zxeTaCFas8rRPQQ/kPlAfwbZ44QZ9QO/tQWQX
ChtUhhPOuGbdGzj9wgXtyfOZ/l1KHDnf97Wb6HmA92aiAswg0Q8Mc/E7lao4Amy3SZJPhNzp3SKT
aOxN8Zl0EN54G0hvpJ3jQC3hTn7qdtoi8DS8WYP673YavPfeDUWeJLD1ufaR9t/u4qIK/dN9O7kF
Xg+oBXOgs88H8103x5ZVbUdiA2xF4yREqvvMIoN7PssEHaXDa/0akDWeQjfaXEBiWxMyWtL5KmDw
RFANcshRJRW5oPX340HticOMS0/bCZqxHCNMQy9FVEOA7jdUBY5XcCDpMzDcyenbgK6Dc2a+SdWV
3zavP3CqLmXwxu6P2bh+ZNBQlHCkqW3ZaGx5CKTDbKy/b/bcDHyWi16Is0u16Te2Ts/4fGWUC12y
gfbO5x4rVA7RFTYDr2pwI10tSRNq8sLgDqRafaDBWHWzX+5FLsR9Qac71siwnv9Cot9k6DxC2NeU
NA9CF+qxvrRidcTreTUIm7GeSvd7IFh8d+VmZyYpWwVkEgsyvsC0yDRiE+ICHvalKGUUVuJNGLA3
DWc8r9qqxtwesHpYDqPq3Gdmu1jFsDXBKzb/5rIzfqahUoVNZdMY9RDvMNU3fbEkX9gjpm0zCbCe
tLO5T335D3SMoxgwEtMlXvb4xv9gtJfuvMtr2B2UcM8a38EJRTdH743VS51QhSM0B9+2aqJ53W3A
Yq8VuA1svSZv09LG3oqObad0U5jK4ifkEXj79VJmgft3w6aphyij4l0HoJRcT32rV1EkKv6R8XQe
UtxdoEfPHrSAceK0Jz2Ayh3ubkR79FBfy25JUoOa16eRKrQnp3FI9yFgd0zOzg8NLaES0TikAA2P
kkXzc3kLluVblUkrncCkWk4lQ700kNhRy5aSLFf618JhAugpbntzS1PvkzNcYeRKqh9eZxK00pJL
y1PrHuqDrgVN+84fBl5WeduyvA0L1Z0vqQcNj4HEQU1EtiVt4ViD5ZPl8wSQsXu3up88OdSwg5Qi
iaeg60ys8Ym3qPjzg+QJbSFVxvg0E1xGLPrb0erDpDMAX1oCaug9PXVGINDCUskdCi9uupUCP1pJ
NPHAvNf7q+Ph/vUvhZrnFhhFPy4RQgncqyE7fN4YTX1Ed3XTGxyDgpnn7BMQDZgVyLOfCZyTrnwY
QKM2L+uMdyLmuciClL250dw9d349YdsIh09BRvOmMvFGTGgsPDg2iMTwZKCRec0NA7OAljjmbenf
lj3LrbqbESQVgih3d3sbMRQ2GH6pwHUBiybv6bdSafQTvJupmb+smvmIkC7rxo511YVXpSIe27ww
KwUJg3UkFYY/RwlGMBDzOuzx6cvCGj/wbvX4gsEigd2Ohqrx3xj1z1wrYMZAsIi0dI+iqrZhr3N7
CHcO+2zk9cwSACSTKSs5B72slthfT2gdh1aW8mCJqqb9Ecl59jpqQfZlXfK//bpZG+KG6v+X3QZK
3U3nroiZMElpsunfnDozkY2zN3d6vQRoj8vkuut0LO7w7OljeXVsnV6yOvoU2y/YBoBIkQM/OJ2F
JH4QFc9TORuMWrZkToHtK/lj4VrppGKHrF5lplPwHnVMrhtu4abYRcR+p0q5SoshsEHHhohXTbAO
PWAWbDLpQCkKKvTyHz5NNba6eYCxJ7KKOAd4BJUvCnk8cUsf+V2dBiA65lHRY85bN2xFFa8XZ3VN
XLHnNHatVDz0IyBCkyIxzvaS8ti3ssfune65Q8jrA/3o2KGbLWJQjl5wDNTgfCmrg2YuOzYqH47M
dyQR18IsD9M3aD/lGr9rQFGQDtphdH4NGY165dmYteGNxkpei3DWLSdP3JqZWAVvdr7h6hvqWtsF
Hgl73yMnRen2MWw4wVWimKhnvv51EQ6/4olrXjvrcCoOIucPiB5g+14yG0PLA28s4zVXjq4g+Fm8
UCcj9VGQ0fQ12zGLdSeurDS8fkDfNXALXtkmHCCVdsHLTsgdotthdKk3capu3A0NQz5wkCxSZNwh
FBQiHy6ipSfXLorNsqw8gBhoZenfP5lrs0RSxyd6gBjgS3yEDazhd9ECCDqS9qwyOy8IIaVru0bH
+hGELGCFwicO3AMRNMzWRwCPk71XOoVK5q+740KslV52H+dJ+7ju5h0ULLq33wi+8GVqLCo1PMlE
8FJy3jN+QrbDGrLv8J3l55a31XRhXqe7wRhpMAHvh3jrhFqth7zhoIOR4yL1nbLga4E1ydqc8Gqh
3uh/MrScyLmeMHoUz2C/1wm73ZgNHlB1mm5OZ3xtqW4WctYWzGvxcNBYD1kcl69pNOYgPVK7RLXx
N2telL2PhKmpwLL6cb7FYSk7MD+wYIZreGz5DcWEsvSdo3UDXrpoiGW8kDQW6QcDx6DfXYz0wx8/
/ugTyFuynvug3+9HrCGxEf0XykGjvbs1bpCW7B6pVmJQZvlNBvbKkclWPBRkkF+/h4ijMpiOdhZZ
kvDM13o4wxpWuvHjm0bgRdi916jZ37FYEJjPKzoPQ4jrS+KFI3RJuRxiA7oxZDO/IthBh70k5fKk
QVRzP0Ze7e71XaJnCagA+eEDkb/Jwm3cUh6/vfsxCbxSo+O8+ZYITNcRphg7PGF0snfsna0hM9wR
56Uab3vs+k3/hEOvNtND/5OLiEJlWNETFYyrb21HnpEorv4GuQjAi68bhM4AWLYNC6yKAY4Mg9mB
cAJkgBOwuXEe2JE7DVvS1Y8FUvDE0cNIQgXVgVJVpB/jFRbS7D+REZ+cJjFrKlwBRcRv/fLCbgWR
QU21YT10cukB2xSnCdSr6K5mAxyHwmEZ7BtuAdweC0jRQ9NuFLh8DCWY9W0w1xAykZZRM4+65N6e
Zqj77GXgINMihYEzGHjNV/YVWPhC+HkoDGn8nS3BpZNkJ8ybWXeQ4CnZBXls8gZ7JlcNU22In+4c
+nY6ZR57TltwnvtKK1s4p2nRNcXYyRUrzmnBA2y0gXxXdeye949TO5rFSCAWWRq0E8OQwFxqiMBI
jzqs+TUGmMhX2hdB4fDu7vISvFCqMaeozjBPgyNe5hsIxBNj74SwHxvNKBAwUs02lpjC+eDn7Y+v
iYuo2mKoR4cdn1ZbLJTGyUidbdb+bZ8crY7rz9h92btRvRDAoIrqaVj5iXk9J/ZBMz1VKT6fJ4W0
1cSVJKOfZlSDrfnSSlWFk0cbHvxAW0NoIcxugqRsjjRsdg2caA3kvlC00X7NFwG7VColHjvZODqQ
3U1HtfCTkU3YuLkNMO4QO7rvq26e54Ae8GaMCI6B5kwRr5YjneTISmpKDVgyGfLI0O9sGJZipD8h
RQJGVFnGCq4963x4AVMQ/v1hZn3V8o4u3OjoIqZjOm2cjyZ7UeDy3DPxSuCpf/3CjYuV4zfUzD9Z
QPcma1ZQgmDGIstmMlGtxlF8OFQz73Od13TJsHd8SB3t7NicTTrmapO887dDK4MbxDt5VDOH2w4S
NHq0FIhm4nbPLuU5juAokewzQiwfojChwTsdwpyvz3rIg5X9Dx7RG5arrolrjU03QYK1LLLNg/S4
i33Un6NzBhXu9Bvq+q1D4DQgZHVsdUQFXg/20mvoamQR7ArpCMnVGvZPQH79RqtEn9w+y7IEU+Xt
UAo45d/Ap82kwgFquWp7X38bW44eemd5CJF30ocvOEC+DKG8CprTC6Bvz+P5a+cn4gaj4IU/yoUE
FVi8H05heZFYI/KGZ0SO6JTAE2En8nTdjcjZWpfu5SDjbIF0for942k7OOpsbRrd3kC/mpIFrhiA
3j+O+WP7DrRvhj2PTtkjWT9NOQtcSvTX+wPYOErixa42n9gkAFXrHVv4npG0yQKGA18nL4GENH33
zHablqikyeNx8BRcz/Hu8E5AGkg21kB2uz/LNGzanLMihwDUJ+jrsr+oo4ZMKF7j2HyYEHK90Wzc
/XUG+4KzP9xKxiAfIXI95uoCg4cGEUtwX8QG8zURGraeUq0+XoBum1w2gnm6NSxoiiGT1jPCostu
h0Skzvx0uAjnMXw6D3jWwiT+U0NiMu3CR5z9WPaSjkhFKcPYzJqRSCsTBoYixPaVCvHOl3ulg1/v
tUbL+KPfDTMEzZ40ajFPRPum8yTWv+1ZHtrNFKXI60ObX5TL/NfssL4jQZ78/4Yp2R6iTzdW91DL
tPOhD9n1qlsK+qtITnpkXdguoA1PF0RsFS9OmBxQogq3uqbH3gSEsfLW35KKQm2VZh+zhIl4eOd9
dZPfiv+EruX0E91cC0+5xWfLhNuKG6ySYHdk6wzvroVjGQk28bgVSl7gsDCSqGKSeyoDF6iVnPRu
TSYslod9R+feMXhG0E51ZhL5BFL2hsw9xCdsqXcfT5PY15hLzwem+i8iHivVlMVdMFxDLXtXj4fF
ldApOXljntzwqbLukRz1qDbZSu1emgjEGGBElkWaIiXCn9If69hLrin3upV+xtZbAZRAnhbZ/uD8
/F6jGZYbEFTbkDcEyMRbmMCHWaVOjyVIjuTKQeN7xWomoM10TA5ERUtMGJJdaUSB1VGeN1z9XyF5
8olGsvl/pLISMNKn1Opd0hry6iCYkminYbfmUoWeM6qEJeKRZPnimguDvaU14cZq/ZqSH3w3XPiH
MmiQss/V9smWAv/pB/8FZGw4X0YVmY5tXO+kd5Iirog8JQXM6dTyHivm6k9z30cE79UsDCtqBUNO
0SxNLOUwUpVFNWvVTt0mprFy1fN6+nvXRMa0JqguO50Sr//t0lniiSW0IJs/EDCx5zAYm7z4OyF4
0J/FX+FXHiKEv73cv44K4j1viyUUpJ7kMju3U6YeBTRcPKth+W5QtBq9Rq0HIqvrO8rgMsVY9mJH
p+fVrHVvAk6VnIo8730N4g/43IQGo1wlLP9oXGNx5JoWbOGWrTAObSoz+oPH4x+IOKTQiRGpxnK8
H6vzPqLFY57kbFo4Tzs9Lr/S8SFCAfg3repCLMN3MY2w4G0mht4a6pX3DVY/iV+OpRk4rlEzYyia
LYs6xo/4DTqB/lH/yTTV14R1mX4TgjeORdNxvJaXIzqLQZN9qAIqKE/EC3+rrpTYOQ8UJUEtTpR2
xGgNTru9b/Wqo6x+XscSAyjA3UciYvAyJrO49bLu03PRYn5dOT0w9xpx3kKqFqaBIHDzMinRJjjm
jhf/LgiwohxPk2RzqSB6qDdTUVgExo1CiYOCnG5KiBM3Z9rVcMPpM76gq8bWPvRYyZCSnkXhz2eP
2tVqP0QlU/QqxIRuDRMwC+DZHYZviVTAvFV7BN3/RyLGzICcjwzO5sZBCfOOSo1bTNHXm8BIo3f5
Yw17eUtTILNn5NO0+xeZcYqoYwFrDbPe2gb8TEjZsMnbk5t4zuBPTs7s/VPjnfEofpRjVfFNX8zB
RJxcuoB1U/tZfiep6fdV5br7Jp3za1Y7OWybgF5+cab48oY5tJ4tZdJ93/EypCWBOZq3xCLI0OuB
TovlKch/g2wMd7OwiwA3haDEEV9HELlG8xupl99YMWzNJpe9OfM5Bk6ozzAMkjONqM0ud8WuNVZa
zdwTJcATf5ZOgMy+1tY5bPvqEnFbngT5HmmJKfGSwrf7Z+si3+l9TOXQiCisnWlrIX24eGS4DKKW
nMYzKfoH1bmW/O+DoUgIWLFYarFCqxLeGRvGTybgLngu4yhPPv2X9EzN//v/jKMljX6iAGSV6UCG
ql9lHETZg1qSOVWUm9AIGWDikbuWJs3WQA8k4UeObnz1yISJu0bmFWEKKHj6ZXiW7Cs1S/a0grW/
Y5JdY4FKs2rcFNWFOeHUKs/kSb0Q56N7Lc7ntWmsuYSg6bWdsTC1sZb7pS55uvSKAuH/H+/IzJHR
lZd8gsNRvdEQG3aZ3lMnJaiop2RH/vYg4QxHaMNdL98IJtS2xXn/q63wI4SiQsBTF57ZqeKd2rFZ
S7GOpG1t6QWZ0zB51i/fq5/ogsh04kzxpn/J9moO7AeFpzB1WKNj/VidWHNOXglMgbJvnIIWflBS
2ZznJ+fNl4RlA/byzDBAkBKGwbM/D9y5XhNzOE0uEcwmDRbEycyian9qtnnNuZihZaH4rTxDdrpT
sPjZBX+gCH5fkTleEY5M4RsCtbte74tC/3npDoVqaYYY5hcIBblqU+wUYsegIMwWKce1vAL6VUs5
6V7ehlBQR18+utl1I+7huCfr3Gf7aTI46qX5y+988D84YraKaakSRg76VIaTcErAbNG8MtwSy5ck
nOiB3ZbXKLMjJwiZxsdtGC5PjueV9dPvXtgEWT7+d3yIAUwavuyBdgBDSsQkXAod3JX8wz2fBJRq
lOq696IKn/1BsBzisvEfWXvP/hnN2aAwtk1VE2LZkniC69O6MKc9nYAEutOdtpBTwB9MN0yvpR4n
ld0p9z9EKPW2bKtmK0ECcBYDgrMM2m0f9YoA9k89dV81fQy8CL+CfpP3m08sRtcYyFjS6F3vmHni
tKM0ed8Mp8R3LCZgQ6fsE5+G6p4KhYxsgyxmv+ac699EobJf+5kjcJDsJcUTw5DWOwsG6DA9SwAP
ZNeDiBfIKUFGtbI6B5qeCmpG3KAj+ZOTFIxsWeFe1aHPROHsuPh0tKyuNa2PvgyNLh6Cf8GL7nk+
0mSEmH4aDvEIVkbCfFuTdcKYXKBOpY/5YPEKTy59wrMJM4b0414gudWREkuYXMbiBRFJBZcVUM20
7vE81z7/nGK8OcuoyvZXbkzhBMtg/KlX0hnsX99jIg4eiY4SN1M2QadD4m2ZQZEQth/9TA3lP95l
IWy707VIZEXNHrSzXao73UPVm2VKWO2UF+n48yDwocTarciB4oMz2XVLaM6kIQG9g+kS3+0bfK6P
0XMo/dLzySJ4CajWzPRj2k3BF7im9lBOsnza60dC4ZAtViPFzrd+Qz6RAhInDDhuF+W+VvenpctZ
l760sVXFv6OxM/0CWFGfrToVIW3r4tTqjpr+K4QwnprD6rSQOucaTDzB7ZQ1xR6du8jAim0YuvMF
4i72Cl9wAFijc83UzkuP3ALEGmaQvjEKA/fCpjroMUmDyNiLnDCy05MmToY1B6M8TkYCn19vuVpM
zjwZIWif6vQDRBLJ8xA/luWrc/yY3SdUqZU9+qo9mZ7W4f7fki6yS9uMNwrVNnqXXbw7fob1+1I4
DaJ63Om8POJR9HMB8V9j4940nu+QsORBzf9MyFqthW2VNj9GU4oF5kL2hdAmZ/ZKJuBjEMPSUz1R
NJGQqUh8C6JoDCNbluwEtivyzsdReBBPN8b7FfDYgM4TvgpwziCd8+P0nufItHQUDUvUgm1Xc/A1
QWuG8XgB9F92qKGoY0puACtGxZj8qNYYbon/l7kqNuD3C8mTYJ6CkjAre9sRvcEe9n9PFCb6wGzw
snkRaSoKIwC5/lF5+/0AkybGI3AcOftU0Ep4Zhq825B3NocSLa99gc/rEKV3lDE73dHMCR04+rg+
BcOnWIKGbifU3TQoL+AG6W1QPeZZoy+n5NwLnSR70yVC3AbcXImfLHV61EjOUeMwMtpinbuyCalO
07Qv0wmId4/Ozf1BbdfjwcDQCvRvz8OZbXPcT0PTGASbADAdspSfjfJGe/VabQDTaA1RnRVuwcov
bpm/2dsDDwBFcQHx51EdrKEkDzK4P6/p4cpuX4UVfe7j9+5PrFaFL1AkoQktUieFQXPkprAelBIy
uD75mYamdu4IC5bwmlVx3fgejM6S1Aogn8sjSdvVndRRlRzvM2EWPZrJBxbzNlj3+Cqm4hG8g9ik
ord8LWVQgbkNBAxiym/YobbYFa4m2r2H0qA8SYXhjmT9eyGQNGsmaDT5X941im/cggFBsHhjCqHj
djCRtVxB2WozU4BTgX2YM4R99c0Q2z2+IYyLpBQ4wvuVNI47lpI9ihBzfag92wp288ql09k6DNqw
/GW0NWb5yHl4pKrR+VVht1fL3TmJdibRgCQ+qGyN4gyI5tdeK6aGzBQScKP3kx4qHhECvP3k3bo5
vOuPOkc3maAQX58YpnLdkwUr/DrQakWQs0GcJFT8izhI/Jz601yBrvmwGporqcT8mp08Ni294kt/
Q6jHvQ1dGmVo3rW1Xl8J2wIq2hfF1y/hTxNysJxIfO2tum/A2x2WToToka0nqigqarK8yvEWd/x+
3tPyLh+H6Sk3CqJaTtIzWen49Eudj58ByBFWdZGNdA5+uEOyHgs6Wto113iPSeEscuDl7R5IIvbG
/OmSkm72klrzuyqc3+2pM8l7NfgrfQa8URubg9dDqQgav83L/yoU2oGPgdOU06g2NoY9vE8h0SfV
tJYOfRzMQiUGo1fT3LiDpaBpiFDk0tRi60H+KU3PwLljHirVmolDQdidbpLx+LUPbaRequT3T5rO
YWR/qTHEZOZ00wSSrNIihrbG5sxMnwOob9qfkjKRoXFx68mSmDwxSzeAw1NY4e+WoOyQZvc8ZmI/
hPtfK7GO2cpLfHSDV7SUvkGVXTzgkEDq2bfQqQdPJWUn20epYaRa9xmqgCCRS+mXq/rTNyYnyBgz
XQiyzYqbVm6QeNkAz0ZdzsP8DsxJetrClblDCVc/qd1JxdD2RuCCl81lzPh2tEkQMnA5lCnMB4hp
7lNbQjddir4hCTe8u34NhVym2o/ljvDHmToIFQhD7pr9ws19Ip12HvPFW4wCWTIFNvZvtZEycF8h
mNPyPm5mZCcmH4pNp58Yd9K8rIR84EOP0UWxde52NTo0333R5s7IRlphIA/ziEGkkUmhOyerXn9e
Ckbrcz/WSsaP6C9z0aQDbLId76jhYivcEySDdGclcoi7l/qCBgVJWQZR1kGef8LM/KjMfjtzrY6e
zGnrhXbFs993XrkXsQRn6IlS4D+yf3a+UqC796DYEaqHWbLbKxRkdmpHVwPGxMGPSg96HdG6grzZ
xyKHTGsROpjcVkH6GU98GfyKXMRtzkLPVSfZ2ryqvJYY7F8IJTvL+Pp9HX7YnbVBTRRQQjLT1LcD
tmPz17YdnHNU466RUkKorVjkc5+FszgkvTExaGYft/FmF6ywCjinyA/5cI70wDirtz+sR5M9IbE7
/EuAqt2iuWg91/gqaUOcDrVKkHcxesMiyJkkSwdiK2OzsKwta/vS3l6DE2J6/WlKP4ZH0aJiUf0y
RfBqlSPKnimX+cdJgeHxUHEHYXqJb4KnEuuJeptf3GfPKdQ+9zPpmpmZH/JqnujMtpJOOC8lPBk4
k3i4w48ZiCTDu+txtbLyyRCTxxf3f+NY+HW9LtdjhM7s4MpTNUYGh9NlQ6UiTn3h6+afOFipMhFN
3oK05UpDSs/ELhi1os1urF1HkHoqekREQS7/B9dxAEPfLWJO5JGw/mbbPb5lC2Lvn1kx7y4M6RFu
O5ARXgP6DajDTYF4+hGNoEZrRifD+DSBAnTAhAenOPaA0vu1aVFXzNbmbIsGgtu6TerBEixvRTXj
dV/3dUs2XyG1mqMQiEEuOvXSNU6xRNlNEv5mskrVjnvxkKFseBC34UAsKxfqGtTuU25eBcu9aW6h
ECDTIo1hvEYnrXZZgSgNiDl5/KwdbnCPpAOXugfzfxcS2Mv6cyTHmKUFQgglit/mzuzkg5cMU6XG
0PkvQ7YqntfpHh4s4S9+8wa0VfRE8PAlFGekhNaJqkXu3CKfwON28c65o+KAeiWkfx01VBiem+aA
YgmKQ4k+pkLYAly9WH7y19aCw0Weczm+1WTnj5uEdIvjUn5n3llx0lXVkvoZ9uxw95J1l+kVU7AC
ksOPym5umd/D4vl8DWG9s2QGWzR6dj4Xsx52y/IwDiQHZ+B/wDojnasXt7BlRC+zpWdywbrZ6Puz
WA4DdeyHw6h5JyQ0jZv/rfXNSmeBqKZG/jAZ0n+R5X5DfjVfXaS7dCm9EHsZ64dFAfvenbWPS4Fg
cNiOaPygWRKtXziCLg0mDslFDPrVPnmE0hUzU6HIyWbgEhmyW9VbNXq8++7eghKYR4ODp3UdJH/V
zx1m0GXHCOW6K5/p1//ymwDHnzQoTNy/8jRtPDPk9o4QcRrJZl69Fq089L4/II7A+WB5gm/vwXHx
nvDaawP2IUVijdusMcJw4QGv+u7xDV2Ua+W0dYIBbnWfEj8VkfHl90/GrT2gIS7g0Ok+ElFRV1jL
UjVqdHH0P68yngMdFVBLXURHN9tSJRaHyrQvBQhsLvnSdugKc/qlbOGnXuVUeigw+BDhGjqGYu52
8+a+XWGTRuqHe5LAyV0X5bZc0nPFWrbCOVaV4W0wgLfaHBMNnw2F6/t5SVg+YLTXRfNcc+cWFv4V
+76hzqcv6397UlpN2t3jPiFoCcfELHkY/wyBSpc55D/xzkVzqQkQEwy7Ith3FnQxoOsS9tqZlHfO
cMXLNomhXuj6TKaJnW8zXDksSUC6RzeZsi3t37CgXCH8B4ytR1hkhp3GKTd64c1tsEEY1GxaA050
QNBYfLVDWYEz8KrbH5EMhp6VL0q0pSVnlLy/0K4z6l9eJi2Bo1y84ukiuWfMQnZtACiZLTq54PHW
TGW92LWfZRPwsplxWwJ7pqNbSd5wRAvnU0O/+rxWaKgxQrAV2DG/0pQ4bC5wdO3kWkOmjFjTwzbC
0liaV7QoBDhizVen9EBlwt0fRqR9QguUXdC+5j6fFaOJM9KfFG6vBFqMU4KW6mGfG82ud9mJOM9M
veyGmEavQlv3ItWyxcAlxPC1dZrXefSLJbbxR+pt5HPwdtOVJfCwcKWQZQOuipMcWphzln00CHsS
pDAZ55I8vzSNkOdlH231YFZyDV7N/DMguieU8TecpZeUlEUiM9WMKACD1p0yFDNQatZ2/4vu3D4a
W90Ts4F7SkwMyEgJShoPd9TLeZBoH38aSoKQfwZEjI4aFCZxIfDZwSOVp+v8NNFcYSqpcTaTnjl+
dudaEpRdorj2FG8gbnzyh4LpyrbtzOLaK/+Z7nH9B0bG5o6bs2b7hsMfh2Chsz5jQJfiyZXV6OMd
Ki/IXr6KBtoD74t80+HOPR9BVjYlL3tNZrr6nMlpnWINpRjw/xhxY1D3V5ICi/F7Fksb2glqpcxF
FkDmVrFhagxvxreVtaoRkaPZ7ERHT7J09kJZXqmy6X2qH6av4y7S0srku83/rHenWhzYTaIvbPAY
LQ/UjtJlMwj3P1EWSE3Mx+rzaOaBXsLyRZzbv3X3sVSl5afM6fDeY4KXG6BhVJp8dUA+7WZH39EJ
WXaHGwrBRbNW3PmRUv4IjZHzeDazZKMwarMCsfS+BzwQDMs5hAe7xbPnSXdwHIZCIkFghMldERlg
BLWF3hOxdWt57573+06FkezONl/lYC2w7TFOo0xqLPXg59416w1hmtrh2WEFGCjrq80m0YklaWyc
C2jm3wmnLhjNUCPAyTGYM553o3w3JGouRW42V0cGJTw8Siaqgq+C4VFoNS1wxPsrkZVbMX08UB6e
P5BQ5JBrwFYP5MyJZfnjR42i3dsWTp8nTSRSil8ZKot/FnUakWVIit6JeGpTA7df86/tcHH/Aiec
Xj5sleudzCFHc6EdqdI3JAKfq/vd8TdxzCSd67OQm1SuwsX7IjSEL8zyliNHYZ2/9YQXg8cyQI+i
3vlntf169DTuD8t09HmRbni/YCaL9JkiB+L+MCzSdoomgFWqYcXxUJFG/Z4fPPn2LUUqgh+R9iqW
eaEkM8FQLNofB2toveGsCe/RA6tc3jkta9kUJGDifTb/muzGvpfKtdwIDEniUZk/WypaI2Z/XxWo
kRmPJ9SGfWbAP+DYYsV7pGzg4Iz6tIGZLBG7/Bdpm51UQnlzxnZc4jMdpRTM3htDp1kEXK5HgjP9
uKozUPTJMBrpSbHkf6iHy7KzbJSz+mOlTKGENHb1x3GWTe62USnZeOZ9zXOpn6vQ7l7f5W/9PxR9
Y8lz6n6BJwaC35UIuzU0YL0LOc2WLSke0edqspc2LDi8MSInZemHhXDqekAy3nTNyp89zKA15EYl
z+VLHqWAHlAUbmxYunDHOY/mxOzHq15s0rGT9/OOKcAsznUNx1yXJrN5WqDQ6TrXIoluSVRvmrJw
nVRtGKr5M/Gq++e6pYsBhna0ZWS+KiAdRwLR5S9CrubAiDKassO+dzFABVuvq9zeI2PRutz5+7N3
cUfNfq4PSA9/r65WDIdAwzAr5+F9U8+eHHJxFf/m7ueCB4s5RGmQAnzGiQZ0hAK/rkbJm7vLzImy
L0oOHKbbEx11Z5Fy7W4Myng1pGhrCMrCJym1gDiUvl+Onax+SGs+1+tUCscQywAUf1U7xcXE2fva
4b6JM+3NODxd3dP9+oL6sCTmVIwtULTeOQvl+3TxHO9oIkvNTASH5pvGJqIT/R7nchcSKGWrBYX5
ax2IoIjltT1NruTKbBjcBFv5o9gaIkMw+KCvQ5DcXHvoUQAa/vrqtwSlfu2WMQLmQIRDW0XDGJra
fGoY277/fSXHKSW9qRu8ypoBOxL/uSbEs6BGXLrRb/MPFmvDqM3UvfNDIM2gZHxp5p7/hYvM/KX6
3OD2VQxJYsf18AUUUb9zB0g4UawXFU/+H8uOA9d0os13Hh46Z0Bcnww+i3xje/lcoQ9lzdt7Yu2/
94DIjTiPaPbGfH+/Pbe77Ge7e0Blr1ZjlyKuGZ7ZbDkosy2LvMQuPnOMGXL9eLFgz1/QpgSgKl2q
EzA+ey6tM5EihrFDTpf4JQw39TrE73ZiljAOWLnMMULFW8UHsEA4rl3z8Fc35Q72caBRCYYozSkf
Q+aUZT4VEhxjkZAWzls/2wT3kzPoDgGB+lWMyD7/C/QjfFZY+xbHXCcPq3Y04KnbpnGOD7XbrQps
Q+mizqeGCn0IenqTFEcb44C2sA9vpyNenq1IDTja/C0RLlWO1wXfo8m+JLYW/OBGF7eRWsPyW9qy
RyOPBxZXEcP8p8Gycx7Z5Ww6JVXwILXRapwXWejqwbTWhxQSIRL+Aeqq+GLErnALO08/83EvMcfI
SelSOR5ChPStFqxOP63ctENsDLcwt/TYCwDi93GdF3SYOob/BAO2Uy1dqBdcr9Y1D+LPtwTmPMvp
yGCn4Cm3ve6TYUXwlAxsurSbTAZeoQ3zW+ZXMNrj+AszqQP048WTgfuQDlCMJnsQYZbA63mXZJoq
VRPMl5hvyYeuu8/zQeEVMV14hFNeiOR53jD7ABo1aIeKZpuqy13rMSh3jIquooAHQzxb/UYuWzcB
l3nyQZAUWrAea5wKNSruMAoZ0fOB4DR3si8fs5UCDhNhxBjcPPQeTQLNsYIflIJzozyIbJdXmEbf
fMtMvnTBqOa5p3zC8fcQfXzhjgmBVLvTer/pIW98tSDTIzWeNEKWOLdi8nizq7CcUygqrsyZaAzp
Ahi0o7iNbYHPYemaPzZmmpIXjgvnic6rmWOD5/JDJl4xsGDN+PDAdeoypyloY1DIovUfO9BeFQAZ
htrKOuq1zbYng7pZ1sCfSyAVEhfSPYIGgXk1NAwhYZIl57X8zLuXpNF0eXsg3tOUzenDWhZDHUoF
6bjNs9FqpQqsimmWC/l6JjkdGiiGm1obX5NHvhijaJnNKoSjh0VCZE8k+mA10/IMAjTZb4Zz6AvY
mXNn3mXGfbGoSi+0eLOeiuKzEPt0xl00KsH1XQ/ancxv7W2++1nxWZJF7YUl6qvZfPD/bZEoTR46
g5d7Bf7fAU+3dAqzBRPnyIA4mEOHD2bMN38F97MSWt1ohlOVHNpG+cn5k5/QVtrfvQiBsHdyCo4W
GV5VV+8oXhrapgfU3DpkyS3n065Y/QNKD0Dvk7/elQDcpNFC54sqa5YFCmRMQoCSAfhJWjd9YBM8
itNYbxwdUMh4/ULwztSjIAYx3Txo7podpZCnOXPcdAt8jwrdMdOiybwUjZbW5KergBIIa4q4rBws
vWWuv1LZtm6eVSsUe82NndVqBA77dCnS503S+mNBXL299uxKhvSVq2yyunG6s5XPeNEssoe4ZqqX
R5Y2qL68W8g7oLlJu8bBDY66F1Pr2OM5lxtLMChtoItb5k7dShaGTIbzP5B6QQE90ofjbVKLq/e3
AnJ8bXOabBOyOg68itxbaziG/IVDzSkPETVJScLH9y7BZprHoZgvXiqb+mnq1z/2CwLKEbjOec5w
+dEeiqDErVmsTT3WSE0Nu87YTP0PTZ2YV+eVjRZXk5E8vYP7YdKO9UJUJ5UEl5G3AdI9aD1sl5LI
ZqiUygBQTVVp3ZNs59vQZqh5xMewp2T/2nOCdKhM7SDV2WFg5/QKFuNchZrovo8IoDsC+1HIL8Gj
HHR7y3+kFEVPVSN42i3rnNLmvfucvbR1WuafYfEpeReRx8GnAlCPAW4uwWcXJPQR3/iTeTruyJ7v
yckE56j/AzYx5rYS6uDvzfCclNYNmxq4hpAFllQk6pcYFsCGbuZI3hnTxiei3LGtsGIb3kpObNFq
4EoAaS7Pp/vWlT+6XCSpMd9LY+lDh0CEKhc0zcHBBRDyEPiBKAjj2+HgoAK/nJi5LaOEGTJPD0Ox
z+erls1Vwi8G4wBrKFvanrJ9TnKm+KvuhsaedKJ+eKQxO77mcewQkfh1ajxwCtaOaFRc91Led/yt
TXyrIVO12+f/Gs5Jn8lFSH+7Ik9MQY6R7s4zZiHuN1UQDyLKzlMuENEhyWhaFFT/2jYdef7vXT0y
BgIE2X/Gbt3XtjA38+dj93OKtD78kXWk9ZzEj24zO3w3pIgSNQ9CU/vZUOfRY+QmzejWbPWPx6vF
oM3v4BOU1d3NOOB/xXYv97WKnzqrZDMPEe/CxzcXpVk5fQJA5xmlWn8IprRWMpBOzfDxwH6tTECI
oZgP2y+JRkr6ihPsFWtcV8VbVxcFMz4svyMGxMANae7T2Pi11Yfm4/ep+26E9b0HFkCdBbPxSznv
0ZihJTVJJlrM31oWMpVvg/YNDVwquhJdehi/DKA3B8U5psXWiV0d59b0Ml3oKosKhOX+NUoVSzW/
qqdGVJ+/sllV1HwOlwY3GqT1MaDBw6za2lyxHn92wljQg50CCct7YSX2ZGP7AXCwQyaz6MsnnGrY
v8TIoqBAvvhhpgPcVABVwFUoE/aEZxRGQaEbLzHA1k/RMEpGNwOV9JLL1mLd2mxHkvyMQA+suWYa
sq6EsOBYDUgp2fbJ2K29bxlYB11Vw6IF46ZFV0HBNQ3oSnzZ8XvCLEamokdZBbFdfDwOnY6OrAtC
jdn1f5VAyNvfdiY6CX2gMabZIF8/EMGhVb4SIFVke/l8u+xh/HNlqDcJ+rEsyjpMDuITvpEKwvQe
c4cnaJTibPE9Xm9FBgIwkS5AoDi7z1QHJURUr/Pum2WT/KB3rO6G4t0IjKWyiz97oSbJWJsiiO26
/wzKjlRN/GSdmf9fJFTPTcbvlhSW/oMBSMXtnm2cdkt9AtEwWkIz2i6BLbSBfyugqYX1UJ665+vu
eJnNFLmW81xIwCP8KAY9wQSNyHSF0BMW5rGGjHyjbkH1vM3IgfgWAy2eoSaR/JhV/8pSXHmwoC17
jY0K3a65qetHoUgvlAtTEGnTn/Dojf10XucNv//YUWIOx3QeQillC2AEB2bh/zNkbN1OaQJGrJYr
sP5gb0PzTY8O4zU4MnM0xry2coCYG+6vJrQp5fJNhQe4S/pRDiqlOeGOIKSjYw3aE8yuEbSyLVq0
S7i7iCFg0b06LieiC3Hh7ldAo2PYdH1mltwqwDVRcxxGx+tGxJxl1bs9Y20PykmEOr4ZZV3kRTog
RRoJbgysEbPBeIG+nxfHULLv5gB32pDut0+DeJ/KyUfSPL5rba3728L/sTY70mvpR2nhhboIztkM
BCb/3hkFdmL0YuHEfdcIRyEm9ITrBQvLoeKij6ZZDHLnJ9drNZ6OWq8mt1pc7gS6MKw2xKy5gF4T
bKDb0xYgVmShAXr+kPnQbC9abcksfk12rBVgdHR4a78gw5rVaXWqkiEf412wAn4HbVVIBezageQN
TpeSXhx6dERKEDDj4Zx7nyReT9eDvpijNN7nhOkPGy+CdZY3MDBzhdavJf4qbdC5nB1D1+clfrMC
SDD4Q+Cy1ErRNn5nFs/2d3KK76v1juhxRCVwdy5j10L/ENkQfqlLZdM8HEhW57SSE4xmW+/c3BRx
kKO4dZXMSuITtR9mSFpZQTvg6ukBng23Ong9G1OSZPudTfVAtu4zmGlaHM2DCNzrOne259go4R+M
8YveIyevsQ5x6izfMORyp1OyyV9eaUpOqPEzX1N7G+L8q4REzi3QKyjXa1AvbTtReHPt3w/d59BV
UT5p9nW61Vn3K53Fyn46OLE2HQ1vSZ+NrhaxjkwODeQPoDGN+4p4lQ9T+qDTFN+XP7HnwRiwOzLz
wYhlpR2DMOSZW3zax2ObTbNgrW758QcQgRy2FR8zLFVXhH/FxDxLMOiEToE+KIZVzQzonlg+qy+V
OiZ3mfsnNyVuill+oCFD796SevRzusssfkdjSh3+epY2jRgtJ8kTCIcRjRqBXpC4EYkEK8zc0/5W
VPz8Zh77sJeGGu/RAsBsom2pfrHRQdP+daJuc6c0DX5/2m47qnrtGGz48OPL25ojY2N8/vWhlxBO
J7ip0R5nn0tXuthGI7XAN2bwgIzFNabdpyHgm8RzW1xB3VzT4COt6mWxxjla7r0ot3i+cgxRQl0L
yrKpuigtmjpu5ESk0HwLSMkFo7sOBIUWPwKlqXc2RGUwIEx7nGJRF6rheJYOWvgaw5Tf0CzgltWD
IK4tZ04/y53v/KNgjlQpOKHJdYqt1XZYZOmFkEAGJsPsZfmUh+2lcr60bTD2KlUhFamSUiT5B3FL
QIny43SBneh61zQ1ZM3NYB+BPReccs7XWdXy/d6UEYqEJCJj71VShtpcTblHMemlOWr3V1QpcELo
y0sOPNA14JPQFHcFrzdfpRWNWWsEQ2VurOqNzJ3QSlpVBwYXDjLI0kZSvVUtVCbj/RE23LxLjoNT
DQJIjm+g9pDq0EC+Q9N2a2Upbt5wZSZIWhNsmhbc0lzRgTU/PzQ2gJrvMXoIgtF1jKWqqppB5/M4
Hvcq7bjc/II22xnhC84EEhgKgDmHsgslbpGIfiV+lyasJksf3pgBcYAbsQxcyXvOClN6SH0DKWjJ
UpytgQ7ivk45nSo/UlGNCGvpcm7UpjDPFKkQRdx5PVJdAsLgPCTJrey9oN7qEYIWn5A3SgGzNkEx
jrExI0tllHABMcabVOtJPucZVU39NsIvkz//MA8nkjbaFzgnHkFc9OiGSgHs6lXScnhO7fzcd2X7
0NCZCaEMX4v3BWzooHUkyLzB4nR2izatahI2XujsQUZuKoeoAL7jbbFclQIFOLxVsq2YZexcBCOH
rkjQGAUuAtLC0lKE2/hmrCiYQanhrIlhhCpZJfv6klPt69PUB7+kdN4xSN2HbDDm/mUNxHp08Rfn
UWbd0GtCzKWnHR++3FSfxy958XuzirxPwI8tDjkTG6UDqoeOJjbawfNsDyge+fScIyb+0o0EJtjS
dqRqcujscXK0LeQ9ysN4PPfH9gaZy2+OFlnTqr49OPxm04COLvNg2jJTivU2nM2x0hB+HGUkSHur
8mIyWqHxJqe8DoCdcPHJ6hNDVHF49jvxh3ywnVWpcPQFAFgJAA1NxYvTS6KrCVvOUpGvRn8vPO8D
jINr9gnWIQkb599x4MUWYm+aWn5/G90A+TQ4fob5yvIhlA647yE4j7AO6GDCFCZnI1G472iK2/un
qjxF17LVHcw+Qdzu13/J+SSe5xMUdOdmT61MgpMDYo+2733p6WzxmZPGeauGHkc0yc8Ex7BeGFfx
W6i9ENbluX8YiccH/HjRORpDWOHSv4e5HoxLLSjtHgu9enJsCdStWk+f2EcABADo0LzmpaeO7GKS
qWEQhxmC0OcwlJHPKu8iC8S/msuGMuPNGnlymSaOdk06N8m4UHvk+r61RgIsCZgQ65zIM+DWDYoZ
5Y/a1KYPb0fUygOwDryvsFqhGe8jqN+5PT1PrV0FgL8LGka4OX8yDMqbbShM6grgS6kgdv/notuF
uFud6XEIMEJIR3B+l6CRtUxVG7jH4YL5wfr7ryMutIVnl8PHMHk8x62cOOvv9aiCnflOFru1lVAd
osbXgdtBwncPgto/1FEuhRw2mAVynj7vwF4LfkwnDEx2Gdk0BHOqZIZZDWyEjpDP8isrr4yTwE+S
e8VD3Dn9SGRMftNiaSsB4agXHJUhtz/8ZFuSemX30ZJLtbqTupdGgIrxbAH4lDoQhm9llxpqoM3t
nlKJz0IUepIUi+QCrvr1/S7lidPsqGqEG635qerMJXLO0Q2DZfsII/2D4fgBWHDYSkjTO3XYPXTk
TgvxYCpQ8ImltWT8dVSZTy9qUl2e0cdCunmkKkdA/D9V9Jaze6WDmhxnC+thkUNMB2odHaxBHjnF
kXUKN4JzQIIq2fGOeEcKa4bP5ZDrcHJd7srfCoebuxCYN51+1E4qijz+BOtd75KiJneaoO4fXT2Q
uKsdg93g79EB4atQdgSAqEhh7rzdCodvsl1mSIJK5PHf/tmMXEzoVoTS0xANCGt7RCwL3wnvcw3h
jNfDYP1Ur2jOt2xypuvMwO31EgfvVxAdyTpPNHY12oZuJyPBKfvzO7LP/iOEhOjKnOF87DI85z0y
wYBgh+fWsyhhbR7dtW+8NRqQVnjiLmKVIqLub/vFsWO0bgw99TZB6lKFPtvexcnNI+X2/1/zeaD2
psjP5xZ5vt7Xk9BrPb7TlelbDt/8wJcMtEt+OYzmxK4gxx9VK44J9p4Y2nHXF3mKbLMG0uXstW4U
PYc8VLONLGp+iPeoXjsX7NOEBVUoY+A2zCGLza1jDh0NCTpMXn5a3LDiIq76NvRowEW/j/SlSxB3
850P2UkAVeKDUgiP+5Uv+DjdVuUaMKE0Nbos56St1CRRcDAFga5Aeumf7rmePBXv+CSKmGLfA5Tn
4BDD+wrZ3epvbJjZ/6bzC2Rwup3Wi9fr0VLqqvQ1PaXCNDeWPNSIuu+Shwmx7t1CtQsMIQ4UpyHf
zVcMSExuNkDTzjtmYOJnqTuK/M1zvQg0n1vBVlHoUeRikcCMOYpX+AtCRoQOOWTsC0YnnYBcY++P
EpRF+/2HWcGFq/2gdua4rBTQ0mOdRzT9Iz9LpwOZ7zjQQhc20qdhL/q8bvluVPfTXT3K0ib2yyT4
+PnlqX5mU/ljmsb5VBOq4SDlcHxttYpm9OR52D6ZCkUoUIvqUpuzc7l+wvwnJxawIf1naet0Atkk
Bp5pRWlXBLv5uU26fE88zDGiPZLP5crkHVc69NMHphn39H5oLXiF1/m8Pv32r5D4KgSy5J55T/KU
HrOEuI+1mcjdELpz8fd8Nfp01ZjdQl7WvOrebuOnl5RFXtidjRdjBBXkGLqEsd784NDsyFWvS11q
L5L6r9jXN06KgooR3M+f7ODK9rWO/MHanEvJ9xXUz1E1GolX7DSExrFvgNDxtQAETS2RmqQ0t7xm
36BCq7i4PU8hpTdlCGBnEPdGVLI0kiFN2/RDEE+ViOXuslmFXfYxZkYqEO3E8ipkKDeYcHBCSApD
fLUC9MbIFEoR86SyqnjI/dwf4/reE144IUNWEiIDy0SGRJ0RAQ/xrs46yzkYYGXb65tzqeTwxxEq
1CPiBgIXIvYoDiVQgb5x4JeTfQsdJEI5q+ok6xorUEAPbcn+8Peb02xSn1p5EYX3eKdvjCJfV18L
7LhNsGW2bUmTXmTqHyLpeyKhm1/pYJVq5mxy9cGym0RvtH4MxWaXeQtjbhAtrkqLbJXLO+S48NiI
fzk/qUF9uP6l86hxzRgyHywC6rBGgJ7D4Pd5364tDggUAtuwOIyswhT0dLFDp+R4/TtGh1qZviXi
H7otIwdlLTwoebL9d79N/k0y4hSR+o5S1Fzl5YUQVKd9zd6ihpYi8OF/rC9/yNmTv12QvtQnk4fz
PW9c+RkcMiil2/62jWgWp1jL/w1DCwZQSjTiK7u12oI7Vtc5MAeUrTkIVHEc696oNhfhbuxcWF92
bp6LXpisQ7bwOhs6WDSOefD0M83E7RYkxUHLf3cWlr19brYVxsrGLTwCzRC+LJ2VapvKH3o9fRz/
d5GPa1Jbsw/u34Dj77PO8V0Svz253JIIKCpjb3DriI8ogUFAssjFYy5hXVxKDITd2uCfF5ZmbP0t
KsqQPT05Dzck1oj791LIBdHHAoxZ2IM0H9fIvRvN70xfWf4eOaGhvHyUnTJWwHga6VnD/Vj+y8Yn
GoOFX/68n4Hy7AYidbYYav1rLAOO+DTBDY9i8VkrZQAYev31X2ux3mGMxsG3rIf+N67pJvbecn3s
X11/95yXEJJlgGp5CAePyLFqwLWZccCqGi0vV6/tbae0z2eAtqwNDFI6ejXLZ2pWQo5YGvVAA7WN
Uf3r7TC/guwKo/tTkzZvw1bVkA5vxvLjVl6XfrXoKmzO53HjE0FiXkaIGgp4ASPjU/f7nJZyZ7+i
xPMMS2+n8Qn1RvDHEwdPSgP0SjN7U0+Bd34LRuXUjdsDGOQnrOO5FZPrXgSKhosxYDdANhLtmwGg
rDQF1doDb7NP0Dt9VeplTjuhUN+IEZAwlvXaGsgWkI2Ry8J+te3DWK/saYDi90XIrk8N3FgS3Nh0
5hhnSxJNEQp45KcF9bCBjNpDxO1fBg0eA4QqKaQsbWtH37vIYWFx3kkAlFPRfL3PkzomwGNZKh+E
LtmE8yQigczVLTKF/a+kWW+sDy7jgkfBHBkgFLgJSHWDgE1JD5nPonDFAP9u2koaYpxlsqDaS18U
1jSM5sqHa/IQ1bBY89HCqJUO11kBn3zE9U86lCsFZIm8bTF/lRYoqb39TlQ9uCz5/QNuOfbneyAK
uYvYlIcipUKjswGtOuTwLhqMmuj/mrd74dk9EnMnl9IzfVCQlASAz2Eq3SyRwMhms5IxQJFrzeDH
uAe4gDy8SxYOUTEXaEjBCJLzTdOCvL3SO/Mt5s9qmft/2wLxQ/6kpZoav2vppqX8FCVjngmrPIrn
rKXehBA/BOivXrPezSPpZdtw60tjfFGKee4UZn+U2RHIH4s7fVbm0dmmsgKqQp/oLky3BbYN2m5d
nOYI2fbXpMmqEwOD24I+m6gIuxyPYh33fy9T1v4ujgHYV/oI91EmAlPSRTv+IylYDPpNFoj3xh9A
xqLszN8T6gAzsnyVVHpUE19lQFCAIeohn1B1GU68iyB8Es7E7U0I1BX0q29ZiapGwQXxMHYPIWmY
106HsLV2bmy8zD7eJvAIIqqNNsM9A6S9KuZv7+vA0rEeK7RZOrnumEztdZ6YRHBK0upgfrJuFdwJ
b2gXjrgfJp8l0PLSqt3O5/umPbU88v9ZWghf+R2ZHVmu81Ld8QZzVFVRaftmyrGssN9ceSgTAg69
r9aZTXe5iUSfngpqMZn+iX++IrAlUxv83UbgbVAJqZgxgJFLxCTyuZ894v2p47QYRrJuFue/Erug
n73QJXujS/aw85JX7iDgxK9S4PqLJhibAu3re1a9TizNb2Z52iR9QDVcMIuAQWgd0OeBBib+jWI4
oYWGCtEwIhVKZqp4ZJm9wg1VWBnbn2obdU0Roy55wIaVTtldSdjkLT0wZgCs5q32o/4aXpcW9EMP
LTpim7creFi8HIdQ/pa3YX0xibZRGwLk2lhovnDfTGeNO0Bb/CdduHmUSWIoi3HkR2ZmIFuEpx0s
wjEBO4yd/s5C3b9RAfsXjZgcqmJa8zTkd4W/ISfmxv/62pP+aonHwc/yZrf2aKPrG/URmdXwD5p9
IN3wnuzc6OJbj07zkxgaPkH3RrUv9Ghtd7TWnw7i7K9xcOm6fFxOyOuchx4DIartP3CV3BZQ3CzI
vFOw5d4kgCjnpq/G+i4wD7EKe20shU35IWKnEIWrTs+3JpwfkhUK5VAfegqkP+zLrEC+6ziloxuM
s+aS5KKfTR+L2+oRb2NwmgEb84ZFosCnzrCla+jexWg53+fUlrHhC69bAKASBuH0z8YinXhSJoWb
vmW6WABx0C0w+t1fJaVKxHSQqYiuxvW3+++w/r95d6vAJW0jo0cMwpayFpBALPdOfiL6ErSt5Yhi
zAnCfwkmFz158Og/BDpeLxSU3Zg3enQ8130IAIIfZ07FdB4h88hiWT+lRzNZJGmhyC1rSZwkIEOO
ypidmUn/xPom9VE9CLFG7uQ3aTeoZWxg6ztelAF4ZpsMDhKXrc1m7Gi8rjh40zOFDd7/ajzv6nOE
RGomN/ladNinQP8oLs1uNHhs3SmMP4gFj1TOjMtrGFjOiHnkgPZ6xHolo6PJVgJ4F0BOo6Ig5rZk
cTV+n/2PddQrDg/Jk2yPT75DSUuKGJ/jy7AtTUIy4bLHfaa5L8T//X5B49U8F/JAlEJWMiCDeUWZ
HsROArSt3/8blas0m3ZYSnD0MUZdzeWOo9l3YHfK+iZw4ImrCaX75YvHnKy9+JskG0h0trfmhGt9
O7L7ehqQdRf0sLCH81ZOKaK4sS5oK+rPF7Q0Io6tsojnf16NKjVKdrOEqo6pws2IOioEf4828FIp
oGFsT/V9jYqTBEhueHq8fdPt1duC2sS+89ICX2RFnAt/34zcYCn/LIRLCPeauOU1vwxIaLt/M+tV
2mofUskbs76pftYPbnamoEJNEXL8iP430AuQkBFVQ4RZvY1oLO9SLBc6+NXSBOAyQ8rmqTgg/d6M
Qk69IgYUY4jxlsuP7VfC8zkBdj2tTaSdnf/pzIbyvFJ8WR2PN2KWbvXWmn3Z23UJbnbxq1KrEFFN
MN8IRYIw5NJBKVYhQyUjVxkAkfB3jrRTRxArEozPXi6F+g9ovWwWr2T9kcG/D6ix6hGKqCSe0f8+
n9JfzNiZ03E1UrRBx920Oth+wkGArN2TyesAot2ADv2CjwFCbVjJQAnl3Kcrb8girHSMS4d2qJYn
ZuLylGbGvrVIGNRXVLk+rhhkHecQVQoN2aRYOzckvkRhW2RSDIfFLaV/NK4d6r9wJBKsUjBzwqqf
mDqQOfRHkqHx1ZhF7XSHAmZgO2DMVCGW+EOA36wGyLuRjP/NDgjgjnCP3wOUJHtnLqU63Zri/gRx
cIwDuRpZvqL7nv8AVN1ZFlL6y3BQ5r7hap9hv6UJYbH0J7mYAOMkAJz9nAPm5nODb7tDaBiYzDXR
JQzphUv5NaP5AbHaLRG0B5Qwa0gHYqECmQwW13+ek/tYFbU+2PUeOU+8gDdXOyoMdy1rIW3k5SnL
3nyMHkdmIngDW3s1GTTEny8v3EMXWkaA4jroJKPFLu53BLS4EyS4N+W3g5stueURcaEihJaO5SQb
gVR9AuCYjvtUMlYortNl31K4e06GwmF5vm+KBGIPH0ZZzo5s3dQBy++K9M2dLc5SqCgaD4r8pU/0
rLSLD5rSeOPzoZtzGOme+h7nfHnSef7ju032dp8Wtzea8rviJxlGYCKiSEevkmcRWJJCQ6QT3sG3
Uu8NiGJV94qNfHLwKVJJ3HylvGhHQ/KexEeUGxYfR47gNFcUrpWQ890pfHyBtYCJj89eh3yNdJC5
OXmAVU+N1b696mcv4otw9TehN5ymnNLYViq3WH1cBlu9WREMFhJ8lhvJd+BBh6AUnIw8SIgHs9KK
1I0wmwrkS62CZ8Bfv4s/bh8BQSpDOdgNBACMNdLN8uFC4BMe1PQG385RFSN+o8mQQXJDjtNC6JfA
N55vKCEaRYTn9PD5M3myKWbDOA8j48f+NDIna+S794SIOOtZR8qlEUqBxy02nfkMPOmwy3bQqFEo
x8i/L5Pcza8OY3W/rjHZYhIO3zaZPyczpBWXeOm9m8m6r0qHpoGemkgVO6EMxrkI4oDiMUzmkU8I
QO1UGCV0tIkG9U6kIO8B/s8p+jdTR9Tzuq7dnk2ojSpUUsC77e9VEQJ7eVMipz451pfjp3VmoVZ+
QAaGExAYsKVjl+9dPz1l9JHDxRnNt+aSUbw37kco1i1HgMHzyop43EG2+i4MDAZha6oOus1mv71p
kEKdW5Thr3CAg2jzHZG/SJUVQN08m6FyU3O/meccY9dFpDODRU1NxNX9tNz7o3lZdz8NhKsMswUi
EmlQ9eBjaqDCwqpG1qZhMO80oDGpFf2pcxw9uvdbPndVm/B5kAXf7ZRYLZyF8ajIubxvrYm9iPcA
Zzj3gKM/0piKJf8UCPWZU8a7OfGkKwqSahZqeK+XUGAM8SnYigT/At/0jDoH5xhFbHcBZo/ffL6Q
yS4zhhBnNgymatxMW1HxtVwDrq4f8UIak26EwOmTtsoCCh3izaOBqthb0hQi6riI5J5afido5LXM
kEQALoXaa8LYNY+kGh9wnzfwAJeeW5opoZtj1cGYb4eDWIyro0z8aCDgx8TZNZcTNAiVb6UWdcyA
Ac3YziU0IS6nP+gDzA9zGYN8BXUpK6lo9SJnD5jZzjWZc0SXGtH/NypSv4co7fylyJuxBCGlJKzc
bzEHGQ5QuTKLY2XO5yoGV+BCz0hrZ2IEchrafx56/kfXHyQqZK7pbm21Js4juNNVrWqljayscPrQ
+mPfU49y1IhvP3P4EURCQz00ZgOGLDLVIBkc8cJZYMd17ZxkbxFbNHcne3aKPCoLVDRzzgKW2HIt
FHYX695u2IzFX4HKZOSk41B0R4aMwTf4S0Y3pd1oGCKDwFtKnY5LH0S+NGiSUrSp5PPLo7OPNiUG
oElVnt/gRiCJC9HwyPkF2NCfDbFr7dic1aZ+cGNZf863us+N4sKvdexKDgLgSXTAkbYEjFcTiY9Y
S8GkBQIoMpAQ1DinVr5RiV95nhl/o8xpsANFGvXGDnSLt45VVe40yggdDTxem7qI0Ww+23htbTUV
XD9ib0hAnZXAOZF3jGNSrp2kLt35/Zaw7uZDwwfilQqeuLWxDWTsbpXI9z3SplL/689NbluH04KT
/TxNSAcqSsZBxH2/TBdS1oEtAnk+aFNb7J2JtsFdL8PDJbCB1vaUap+CdxrMiZBB8JD8uCX/0/sw
aI6SLv/qQ5XA7oyEaclddBVc+4O8c9F2jd+TM8pQUDNmiebXjanr1AYNzehnfP8rgSK6zmIdl8ou
uKZwxVnjk9Zj/dOIN+T/82rDMlzUfE/kp0y6tE/xiGAbjYc8YTi+jfjMdkhcHgcdVDcNAI9NeTvp
2a6DlHs7cJ3pLxYRGv//QVIOar4f1wpkh2FfVOfX7OZ3QerLRMunWwxD4Ei2xJRsZNcspFhFdnkF
Cdq4PLKZ7YCuPoVNY70UgB3zOzak5IT5BNmADoUnsMWaIC1U6z18LwdJZmq4ObWP3hyFOeVVvunt
FGeXdgeKPPEJyEyhY7N8/rjirkLl+wp/c1h1Ww5cyyiRf/ynIiUqKG2OISSy5KhMQQxvyTrZA1Zm
ZWSJJmYzY1IYXYy/qamAoJxJM182TpouuoICyUwxTwW4SonPbwaib3PEIvovfj8YfLYCJR6jLVeH
1DdAZ4uwAJhyTcx/vr2VMgpmGt1/vATZdeIhBqwEsNnpea2kKTnjHpD0EqkmPZxytv/M0gGtgieI
qSD+p4/Tta6MXeLql+ZQC90nMK9hgL4t7K8gpb/CwcEPSh39M2qnr4lO1PjJWZLJeYtv1eAOpctO
WivWpgAAb8PYrK2p8ozI2H4BweyHS67ph6oCEXFWr0fA5pzkNSfTEjMpergMP1X/V1fipyW52Chf
g3yAG9z/Xh3VBmaM0mEZtlQMo7JDSxoSm1gB5Ko0SS1Lu1v4gpsF7pSdRAzvZGe3nFgy85rvnLNO
s+chahzJWp2gMYUYGlQ9sw/Qf6OmPnrfGpLRnQ4G8Tdqc5h1lBMlPnE6kS5ewzIoSWPaXHGU5VS3
k/7pvAsSJZXu47Twfqg5+G0LJh/TMGk5KFmbzAWSlrn4oHGqJzCINjMt/y+5zRubAZjLD30uAF1u
GvWzF65t6JKwzMgoox2+2oYPubOhta4kNEcISmhPZJsL9yRG6XWWBRWWQ9qqdoZ1dRmVN8qpCOTe
YA0KdPIFWcloqaXWaVGNi56eN52vWIlRRa7qlL5d/MBYL2uVV+Vu+QHhBjraGhu+gGnSSOrd0Gl2
XYNpamqy8bYiwU7mdMv2r1vKnEocXKa53Rwi8D1oonGom2FNuqcKjmrIE7p2FH1Rw+OJrQiagMhE
aWFhwL0Y1nYhMrcAtGSBUkJzPAiusFX+dwbZzbDMBGQE47qRGpokhQ6HF5yC9rpB3r8W4A+FXq4M
u2Xi6i85Uw4toHWoFNy+pN2It1jjICwztaiCsblmIMZb1lSbodSSIo3qNhxLhQkoRRG7FGuG9OGz
yDkX49YLu8Viwgy3+Iv4JhcPoXnxCsqJKzgSp6gof6QXRz3nxM2GpVsClWM3s+MbE4ErcPeV7BYF
cMBHdJirW5pTSmwQeIX3wPSUbszexv2Uju+YEXmz+0Zq7G6UNVKM85U0OtSG3Fhn2/cvzPYHVNsT
bhRQ0jFd7GEpeGsw/9yTPd5hK/DHCbn1M4asROVz7hctWn4C/rgi1bU9/EoWYsRll2dEMXFylf0r
Zg/G6ms3mlZcIs4ROE1GCqDE9T0O4HyUbULSuYry8F2E1l0N9HDlPJT6Zk8SdZ2EF4NyRAime7qK
VcdhVUai00+3cee/xWYwTYYOiiFxgdwA/ZUpdGH6XPgzeXU89CIZZmix1wrDP4HrmagpUeDVhVPR
TO22FSgMaSItmTmKoNyhLcaxaXsH7g6XUbeTwv7feIghY8gRUfO41bHRC3+gEmD7v5UAPiTOFI0W
u3yuxFZwb3g82DAppfD4dFMgjyibVSVy5UOz5fBpSZOkNf/CTGNJpQRSa/uhG7UCIRwmnJ2wxMqg
IZVDl84kWcu1cOfsp2LhzTpnrGDDvQnQCbcOiyY50dr4OISFOM96wSVLWDMBonnulE3DhOOie+bM
XiBbA9LpMCbLeIeN4UWkqdPZTaH5tZnLA0mTztUu42vWMF389WZNM8aarOtIp5j+o/ybKdMw6PXM
ytC3Sr26Ea6iYkc3Z/dygqpKt3qa13WoIk3cE2DexEYTNqWqfIohZ9omOkn6RUw1i91Ie1sLnUMQ
IOu93HWcqLyl6+vIHfHDX7E9mhYhZlD58hb5h+RlZOUA1VMzVZ6DRnljYbfFLDdtUD18d9jEaD3f
mM7eW1FhIFGFXm6tDwQ0GR89xfz0fzhdGTewgX5VbFfdZaIKyrgPPE+HYebybnyoFckDblRaB6yz
ufAKPbpdTmiattFOqgDCK8lkWLEIw/8DzsqCkwgcIsMIeiPI9Aoy4dtaRUw8F519yn8UkZIh3y3A
kMGiJHFCS5HMKtVivERL16t4B3QF3vRAMHyN3iQe5tKi79cOpDsbuu1Y/+/qQMwtHcrJIuI/xiXq
Ay479twpcXvfjmz5pgRGUN43ZiXPhnXvRPH58fKEn+K6FERUiwRQ9/8+GkyWZPPVRgsrWgPLPDSL
G2j/hJtT432l5+TQ6At8FH587nR2OLeDfg8xL1lU5KubfKXwOW+xR/pnETXebVmXXHLTwZmXsD52
237BwSi3nkJdeRBsJF/q7MqK87C3fQpPHCf40pvPlSYVMkfNX9r4Cn6EOyNpFonDT1f3nqLI9c/a
zDNMJlICMUHwYLC8UDwM6fvS7/8DcHn1Sjmk3Buc3ukzSe049m261eLd+vl78ZsOPbol0BLxRqtV
asCDBiDDtlpac310/RSXEn75PEibBQraCGKovSJGHQnz4O3sOUN9fcvPwjEqw2JNdeHGm7oBOF8D
LKpkYM9faKuZDVTMTawE762SqGvsS4resijEgs0AAefuazam6trY0pADbAqHuofwSYYu1/w4YYoC
nEN0IbfjNKaeSe27J4NOJx3uyAZfszeYZ3CmR2AeoRGrC15ZKNI/XOvTesUh27WbGOuIUSDIlyF5
dpDxzrJSLvJvEnenru1bvTvXdB8106r3ZdfMNudrwvVusEoangC4NTKhUmmFAnFVsPD+hKd8H3p0
OD9FVa0F1BVJZZEEc147y4w0Ch1nRSQ0B+9RJQGCj40lirQnJtTabBH3yDw78fJNtEHDLsifcElJ
+WEm6TGIL470Nh3pslYLnFszMBboJ622DAPUGB6gHL467CwP514NxFQ9YOJQqQAftgm+jsO/HyDh
201rrDa56F32l7mDEcycM3nCc6AUOjsbwpyyBVDJemd2jlER+XdOewpVnvlBrdnPmyMjvtRbwx9s
XRa1eWqeZSvNWVdpvo8P0wTeErDyASH/MpjQDNzUj3AbON4zXUneKyKbhVtjRQFlnnSeyykA4qJC
aPREyOS/uoP9IdESJMfNUTvY7WQ0d6p38gjFJ3G6XNuIPn+Y9PiERMh2lqTvWKdS0EuNgfObejzv
j0wd4+f44+qP77PEpFhpZIkn3F/VeZqcua9dkMXb5piXwAsUPNPBWxg5osTaov5IbEPNmPqTQVDG
i/Wk6IX/nMiRXnQsPGhsRdvbyc5RVwE9Ie+emlYw7Mh8tdYCk0rMmWKUFRKuBa3AeO3QiYwquGNI
V5oeiGaiFT9gE3GNWSvutIjBtsF6oWLyDVzOm/wgsMAr2ruDcigouSgcK8xGZhUOax0rR0Nwto/i
WcgenNMc8rVO17kE5fAH2B8nc5jq972N84HvGIz2ABnEOMFTZ4qtQNOws9jjte7pZdwr4QpKu76Z
STEit9reBsuhg+my3/RinhSXtXTAfw3w75bIEj8Jb86P08OFdbLIe5I5mBIoIlWcrb+3aDPxQQuP
7hOQ5cpeyWrltj13/83TyhsBeWAzGCIqU7NwJYgvanbDm2iFZ1rrxzdu7uQLzrFU4a/QOZGVB2Xd
8w+AhBjt8UIKZjXOACWpxYHTPBQwUE84PfR0Cm5bAk0d6gtcQoNkrZ+Jk2XRDNfM80lUTfBleyD3
yqpjXdF21QPGgo9MkbuDvtdi4A/UJMgS2B+xjINfJftOMNr5U4ojSNmqNYlVf6ZBrxTskbI/sp1a
HIGwCVB+9HOg1WAdineWqGIyrhjtEDJxD3lYrnbcqar6+XWquQYtXc+dWR5x4zDUra/p+AMCno2Y
vU5ORlcl/cX4zTiP6vck+rf5LHw+FNSK/ajY2tLZvOlB3FKPqD2ct7Dsy7aKy3cV5G1Rmx9il+NX
abm3WSvyTOQzsxVWmKpvAKp1XYByNaH0rxvsG0CFoi5ob1Wp8qa9Mdg3MQ8oED06BC78LV0gMlf4
3XiH3a4W+WkH/f2Hc8wwpr0EsacahaI0FtCpHiBiABKRuPi3P2SuDKqTWvhTCwjtPrlYMtxXoqBe
g80Xy9CWdqZ5FnMY5SiIPP/z7K3j02PGQoPhh2B9gsJO3YB5XU/we/N74EiFyAxolUfU49OclVU0
7Pw9kowCMGN/A8AMKHMdjL4ENDgBXF9lA1oCMfy7vBEqKcDfrKvT/6OwHrvTiuCGvyWT5dO0rFlz
06RLM1XDkz9U79L8Bpm8atlbFiKQok10rU9CprAzxsodx70uzkbcgENiv8+brrrFfoJnWxLy+hS+
cGq1dPODj4J+U6gTX4Mc7ZdtEqgfCu1qcDeuca0M/5Fx8X5guhlr2Q9HrT8vFhNCuDMKnSAciSZ9
tZ3MnlsxXYubmGTXJVzRVKBe1fzGgU2711B/5vvdEC5UZCM3c+msRUxXxFMH8nkdP5awnulzCfhu
T6BNpQwOAKltZiSNQkapDZ788XDYlTXWIAx69uKz4iD4dk9YTmA/yovGzAhsh92YST6ppSJyOTBp
PiRJuR6hNCDAxWSrkbAAUXRt7qOw+VUj07WjAphp7Z7YfjjOH4jW/kzjkysKqkV/AluBmd7Hl6vK
l57CYq/1KvErK4h9bWSSNPePrRGYL1cvTEczg4zN5hidQ+sc1yv379METrkOxs3U2yHKK8WUcRIH
12ybVwv/1sPv1pnTbBx5WxRCALK5QQaWxLTikgAnLleHTVTN9HG3ar1AaaI6La5BxCQ0i7ka+UmL
2Hf70tYS5A0VslcBU9Oww5lgfTc+spNsHTrZZSlVlyH7AGeh0IH8C4qHV8erLBTCPDpG+sLeLGLN
IHIgBQZGWWHg0r6gpROetKouKzFqp9bUb5OJEp0NJM7VQs11n+sFWvizgSwiYBIjrtvNflSPTgEn
9NnP5OMtVh7+UGhR+OrrH/MGAYNtMwkH2oEHM7d5CZ6WV+efufqd02ivILoyql3Lpi6nuXG+/Hl0
YIplIElvXNkyJh79nITQyKmnF5faurjms1UeRfStkXBpEya+EERzF36bOb52X5grZ3l6y0KbFRH0
d08NedZ/W5rUILUkXkO5YkGqe684jikQUDbdITerTcJP6uKGnJduz8CI0AtZ2Ubz4BVYiKIkKIdI
VUPft1+fnKY9R0MJzI9BUfca8fhc+a4k/v2ZMrPdwK94RrQKKt8Tv5sv6vfLYHH7AA2nvxBWN0Sc
V9AX+g3XGk0dKYFEwQx8ywS6HdCW/nByfytKTQsxH84nWzt2UX1hOSquVlLbN6DPJ2bYNGR8gO/R
E/m03E6xlGkHrVZ85oZufezELkFboewzOCx3dXdjIagsrflWumQfhxqdBYuRksJ+A+4Uk+OcFKeE
/38msyCGvAo7Xmu+jAOc23GIW5X48/F4KcG827iuI9qEgwGJ5sBm6b5v9a1g+5zY6BE2Qhf4of/8
m8mU98APEUiZLCEBka4yYLg4lWvKdWyEGtxdBCmo8Nh0eMRUrbCY5daoQ81NHcqgBt7U2GLjIY+0
Y0Td9TQe9EM8vaLFnDsgLQy1Gys3VTxqD9YwwoUGKGH8qZZHn0A1tML6PaG0qzGEp40jaAUmnc/Z
HRghmAJ2/nQonnyzJ19YINfzQY7I98ovg5GSj7N/18SqA2eNeBm24l6JQEFkRCgvnHxFyMWTskJ1
CKVEU7YfFzHdasvPp8o7976K8xU4LXK/Nir1gAOjLuZoLh9jHM4IfNfBFYMARBdt0tLWb13LP5Rx
LvIdC5+LRyCM6ShoHWRiz3J52JznWvEtNLWLpBfZJvnGBOS1Hl82hcTgz5jYzQ1KvDWAH+hFE1vW
NH5/pz9wYrzTCNKvMtpsi+u7QudiZTJsS0T6AqR4+oTmI+2L8jXZZkqQOyM8X6wboV3Awz/sxnpJ
GV2N215FqsHZE+OY3WZTae9URyvo7NcI7btfrZzaAXKJPqPKlzXbtiBLT1FkF1fCZrHYVfksv3Ww
k5UrMjgVo0uRq6bmDjTwLhjYkLdP6CruNjsre9fjbO+e8TvfIAppiEyj8HOCZYMKiSkAxp4SHZkD
SDWJnz0pLKbygr/P7Q47GDk2osviN/oMf/l7/Ilyy1cbnbcGYq/udzt8T4TwvwFFUW17xGnwPCgv
q31dqY9CLADNFMgNXq9RBAANeD4GUaA4RqvWPkLj15uy/i5nJ43Jm9uFT1i0aZv9sjiYpMC6b0mX
8EUCaMYfuEIMs8aB8/VYDFsNFAPHdwrQX6oskSB/+EceEcaXPiHlzVseEeTZmvyApZ9EgKon5D/O
LzbeR+CuJPAn734Ehs93i2SsZ1ZaX1eoy3Hj+tgWuAROKh/YcQOJ7dpVYCv6PhUv6w5YFq+GKJEm
jfLPDW8ozSDpkEP4lzj5P3fAK75Ztr5phNgwja4YDjrJIZdrfZn34VAYhPVT04WI9aYnqkeYOPr4
rmGBXyV7agpwLSEJ6S5tPHdbbIT4gKuJoml5TGzG7Pj8ab/mGxlvIKr+tc7AC1EsecXVPt3FgGFr
WheWRRlIviGKNFEUc9brAeYe5SSFyI0gwWtlEM2b4XYyW1Zj+WokWZ454MOquosr69E2TuSLuxo/
iZgr8+cCK+WFox4DVxVjhWB8yBUricoKrHNNUy5ei/CoFsQ+6MMHyW7qTniqY6GwB18wkVxE024b
tV8XTkSNW1LdI+2fhPXl90LGHN+MqVkXPKKOGcimFXY3ixpjZjiRJrE4sr4w+ThIjaBuWtqpxAYq
cBid7AO6a2jKy7RVIVdsZzPpSRY140Zrbsi0vZr9VHbLBRKIh8tNqJ/tP7DgPYw9dX9VeRJy6l3O
H1TPONoz+Q7ugRA8QJRNDbp9PWXcilAa4euRBJFXlf5g/FOaDAuowMaKo6yfhENbVrM9Aq/Sat2M
3joG4qUqulra2PaYGOUdhAw8r3z99GKskajACcJIJrbyYV8Y3Vr00nykmbd2eWQl/Lk1bsqCB/Ao
1SIpAIKRCFP8bAbFHMvprG74xmiXQ8hHdAfICWF1sDKZpiAbCsU4D/Mj1UARO27ywbM2d/oRND9V
bXwG22iHBLEfQB5LEvpCUO7gE8Cr3FshdiZ+T73cVQ/qroVFE6Oe2iNng/pe2oTvxdO7IUjsQTZw
jxVzFDx0ceoq4ISSCTT+cBspHVMT+pdhMn5tURBaBWqCX73cX4vrVwl9FGbeF2StcWkSCTXd5Z/5
Bw16rLUFcqLBvkQn6XYDc7sRekr8PwdqLINxLgEOlLUgugjgxkuQUNl0lXcjYnl0LnxNwWt1fDHB
lHISGos8BAYOuuhZnbGqUSAssWxXucXIMPG3VsNpkqi0jq0HjlGzE9M4uNb0iqYi8rLHicEI3hVB
pYi3YZ9zl6DWexeUkzg9SrTViI9Q+WHB+0CRnB2SXqFv5fCfeayge2rmSlRy096D3mY3X9u6nhLx
okyVWlCnP34MoxTZmegnzLkEzFCldfX7h9VurSdvChyzBDZ20NeKGDwGaCocI0PSxTXX0Rc8OYYd
1Nw4JDu/jPkeiXI89wPYtGq+SWljaYhIVMVMgK2GFwOkb1PaQVXszauByZm7f3Xo+QQhI0jelEKq
ThFdkAxV59MJpwQIzb42KlSnCWPTK82k2P39anuH0JqlDmn4MWRfY4wUzH4sEdwLrlDuHbmFqYvy
/iHtn1YSCYiolbL6Fgljn/LeLQQ9zNU9ojpihGnNGuUyGziTyd+uoSLigmQ09rWCol5uBN6dBaKQ
Va3/c2/XzCW14+PCh/iY3C9/4cT12yPC6gjbQrENW3FnbH440NYfjiHvoRYN1pmNzC54rcYAP2dv
ZTkv9p7M6RVthVnQ33jeL5EF7stjwkqTBqSGC/RkjtvxX1mMD1Rms5TipoO4+Fpv8iJf3MaBV13F
E9SSzBgCQN2EJteWDj3mu6UZTkXAb6A2gJ0ARAli258AKlpSpNvFw556EKpcoyI0ueP4Zmxa1VXK
BExN6qzQ9NqewoBrbEdeQ9yYKqOfuIN49Xq9jxjSBHdv7eUf4f0cOH7whh3/Z4zjRHmEo8fiSs0R
gcLZzWE8ksp0Mzl4rA6fiuNpz5O/E5iM+8XBe7MDLrmB18xusoNjcbbAJXb7u17u0qSI6anWRwxJ
pkiwFXx74jvRDsbbr6FLP76yzpXGqi3/8/097gWbvvWOmxQpvjaDAQpPePfc9aMjqZp4yOIMBnNE
CXCFFNyenhEPILuV2iDs0SkW24tRiHmHBdKSIpnhZxnU2SGrfwSOhxKiz0ZrVzq0wYTNSJ05tkL/
NvnhbBC0pebJ8sD0/dcScJY5U/5iyCRrJvyJVCdGeBsPB6fGUZJMHmCB36gi8zM0c9P2P4jzenzG
njO28MDFlXYhc3KvPRACyP3o69gnKj5pO8BdwqCiWoOCMoSEjByOd617rX6VFiBYrANnhWpedQ6O
DmZAKp01k9PidVDl+Cf1o+u3284VX6w3g5He+NoMD5WSrVUpicGzIqo+pUfGYgVtzCS86d3GqNn7
pNpvul/AsnCXA8qMtm3q86LYi4WH3lrx5YipQRKFq287c60+z/RLv6LSl83MfQ/P2tKj2SgHM2QS
dzucLA4Poh6ARSNFRKfVa8Ewv3h1mwYQB0MHDwgQAOETT2RH124+qIbdNpFBD5vs/Tx2QeNEvnu/
Q9g49QbcU2b24Di+yAkESCNMTPgNk4JQhQyhsZsRpJe6ZH+1iMyCZWKXecixSJZj2XhpqFRk2HtC
G+df3REJd+5jlfaMuyN+qiBpB3INYWbgWK4SJ/mtJUKUiJxajc0h0AYNYcMgJohjrBNnsHKAk1A7
1V87i4NfLrGAH+p7iAoxL4hH6+m6BLgAke2y69E+2GVaDSOSV2I26K5e30W5MvUcaorjKBl27mu+
NgI3VOTq80KV7hdpuLcxynkNwU4sUXTZHiEBs/lRtGyg60iwjC5+Nurli7pYgN5WYylaNR56XJ0O
2daZ1/ZEqMB3f/Ai0ZShJtzklBVRL33zS3zDwAZPaHef/D8vAy/ulffvPaPJhDxr52E+59eP1S4F
oNfm4dX3SP6YaF7iWU40kVxiFB1m3LKW+btyArLeMnvU4gd2rBz9rw3W6qL/iwWRpN0Fa3XP1pGf
205Z2AbHtAH9OIvpHXE3LyebBcmPTLpAz3KsKgbxHXMoNOMJ1lim8ReSBYCS6n/+UqqY37T58nk3
r1Qpny8+wOrYekdkRl2bPUUFjjmiaXJw4/YOobb8ii2K/r33Th05xm47O1/aXLFPjci/1iS8jz4/
rzOF2v/HCkhCBtMA0IHJ0M/By01TQ+SGSL6XToQ/XqvAFxmYqWtWxeqgPv3ZTarT9fIQGQFQLuFZ
WZ1enVmRxGWmPgwJE8iXNNnzDt97Ty3i8BspGUAHLjOtMm5yksFKBgsrafBwfaHLL+exTNGDsjcY
pffPSUnbgheYUtp6PLQbr/xmqSOoqGr7tldd6RUE0jHtoAkkys7733mRNPGLZaIJksgtF+wa2/1t
XyxIw43P2nOlUE9d8AzuBfQA1be27TzE+LBZVM2SP8Xepf5sGtCBHIZDpZw0wE/3EHOr3OdMN15w
gjpyEDcaJV31OcnY8NUiT+7/1Mz2taVEc51y2hzVO3+ME3f8YGA6qoBZ9Fjzwi8olVqHNU92jsJO
3GfcQVyp2TsSvKsz0leGdpr8bH/AVY2wduCPMltD232V7qk7LirE58v7qR8/zF8ZzFYTjQZLqbNX
u+R44l+wH4XiEuzfRF4G5sy/NgYdRJG+X1VkDV8lDIm1o7fldAwy+krn1U9reQyUwrF6ZBFzuWf4
gNkb50CkVrKvjsfLfNfhRKUqIfBrU4NfgFJGsUdvN419ya3atKRxGcuzf9FuCKnqS0NxfY2/+f7W
SZuMdT9UWUtWazxmqv3Jv2VkbbnfLng3s/0ZnNnhuxuLNKno2qKTfkr2EOeLtDw5KdpgMotzPrRE
j+Ao4RBq5s4Kb7VI0vl+ap4PPnxG+IVfRARjVtfJMPu56+KWNqk3MgRE49rOePBQFUsH5kOI8cLU
DG/cq3wFH26AwNv1VLjAd229x7gz+Bopyc6V6iaCCExN5WiwQv2I+Ky28nUsTZVAdxEEYS5SVXOn
3/ok+s08i8fnbZ3tZ0BIgKC6Jfh2DCGm39mJgAKGpDL7eQOskulAxio6o9MfbSfDryKap6RU+IzI
gBLWWS5Ip/Hcn+cbbHK16y+Iwh4YHICs78GSrDDbh25VfcjyAZkvKZUWtPDJB5Hv7yXzhHjnbxmt
BD4JceSkMzCNqki5RG154wyJih6mxj+8ZmA5nOeHjHJf6UWC2zfVBjDZ8H4mtU4+bHyEQFLti1Dt
yYyhdzrD7/pKDBHKFuEtwVj82ouwhjB9Qguh8LQJgCmTHTDRYg77Q1fX4XqN3t0cYtsQaB7Zoc5n
aoLEcP5zGXfPnI5Sldfx7KteQTXMgsUyUII5QMkrhz406qvN2WsVtqum+KEwFlN+3ukLAx/kYqiE
JxFn1LF9Hy2iRU5YNufcRWS3BLyDHrjqiBAH43Lz8AZtqlDNFvDYoGDRFbtLjQjzLiPnH/hd67I1
GMA7jpDEZwtJFgfRQqt21WPMzCngQ3Z8IpfcLP7Vn/8G2dLWXHd6cvGJYbl65cx/KOj67DD8ktJN
HjLKNy0qqQb+7uDw3G8ey+4N0lovx2J3Rc12Jp+h06Nekyeci29/ZtE/vmRHeZmMVPp+/HviLqcC
g+G8gOjb2nYgu/A6ioLOW/pgRiwVlIgmKIbRjParL5jNjmf8PzPi9TfvU4yUSxrQ5rJlhwOchjiY
6D0oO8Ht6uINpubmUFYnby5m2QB2jI1HPNSfWhpaFnCesmSIvIKDxJNdSP7G/KKJIVnTEkGzsx5w
zMuFl6zj3KbEMOFGaSs/KK3az9/8RIIwXhwCbI8dt0EvUFko5TSY3T4BlEr4FI0XRyNJjE+1SX0K
9W41vIo1UP/FHwbWPoehtz/3Wf1wfEEQ7IMdU8sLdlC76uGYOTcfBERE+I6/D8ozh69sqwssBLWw
bUDey5K58krgLzxnyc7aiIOhD+yXJQ+jkvhx0IW7wG6OEZyQ7zgKZg2N/jbRzhrkCt0ya4jRtAS2
Mo2UeKIniojfzu5nyoKB9z2EsccxZoHtw6QwMxQm2pxMTf/Wf1wdkATaOVmFr+Lu3SjZgeUAjRGC
IDkkoiwncCi/2zUJ6/dGCen9Xa3lLndIzAKlKCUuxWG1Ohl4Sq37gD0QWWLN1DgnOQDeCMeV8Fsu
apm+f+uAFKm2atN8Ml3NiKtpSTyRNeE6aTPT9RF+7iEO3GMgPswcYGFK+hF6F6pF1e164MXukVwR
qkjMCVjZbFDKitoakXBL/I/Va85iz9NZtmX00PW5YnBS+8sU9Sv5A67E62ih2VmMJ9DtKw4l+gMa
3yCe3S3Edr/uoKL36VOzgu1PGuF4wamk47XdmpW7vEHQMgTEtSXu5Vya9vVThy9Pl9y4uLJ9gbAJ
GBaH7fqJOKxX/Ggo42o0tRlkhzkUkxI91BYioYswHldTVGHUsLQ8boqL9XV38na78Op1ek1PVbUT
BBs0r9HhmzuMUae3KpzYwrOijh/qsvBdMvYV/ZKc7tnqFC2TFaF6r5UlfD7CYbYg4ABk2vR0aRHk
vvtA4XrW/P0AmqZWrt0PvxJHvN8w+LZnePIZ8dR6ktztDpcHkGmznnZgw7wiXFtO+7g3Ia9IWHHk
pKoT8F3LZHgvdMBgxIQabrHFP2Rl95/5WU92YEyk6mYxuZCultRhMhcCArmsXrirITmW8C8LkTgF
sDryiY9UvREAZeHmN+5uE0SrSUeejwLUsY45QwVZAyNAHt3IEQJdLkaoWFdAW6a/JnOgD4rw6ACk
iLSeuKieqk1fb6v9JiWHwtRRjzx1kRqSLcHdnxWA5BA+bwAOHVhZ2eUvYU2py9bm5FtAvSgw6mNf
Nl8CoeulJOJ/+kOXvKGZ3Ub+bKNYTqMfV90vyoWsvUOzLjc9Xmszg343i4SjR4u7+piuEdReF/l5
tA+BTQDKxBMZ3VOKSmFG/HI3riGJYf3Ask7sKkc9aqksf89pk1zxtXLscjXeL/riesFAJLFy2g/d
y+RbIgl/q7GC41JNMXwi1TmaHQD48B8r3VHT8+JOt4111InSEtPRyD6W6ZhxnCQCvcoCh2NMyMkp
6QYJcu40uJj7hb2Vkg4+ElT3FufPX9bJwKOHjOAPQUFktWFwWWBtUQwyAsstK47sIlKdc2npoz6K
nVRy4utP8IZSiWQUsBWnbwnh+LwkrEseGnK2I9nI4WepJ4eaG/Rhwr5AAt7q0Dyz4rwYaDCnS0Rp
FlLdhBXev+sbhNxDaNKtyzIAP/sIXHaA6IZ4jU0ZCyJVJ8uT3+FK9vYSD3WAPlEmJ0d68b/6D33X
BxiSNHqDRnszNoUNTmUoDMetPnel+mL/4a5i6wTEAISYuvG744KrzUNRj3xIudFEzJsAAXIQK3gS
8iVQt64HSddQFCD0oh8+1DAK7LqHzr3+6yzmRf47oWO154sm2PnoqJVHLjDa3iQukvMnigIRbg4x
kjYZ2h5yiv7dLf+uUdn7TjDsHJnFg+MmBsPJowuIFyl6rIEy4JvwJj3bfsgXibLAkRcFIPlZ0acx
H4I+9rcFW6F7pTQwIocCCw5T6FCVI0BNuiAsW1s4r//bEKeMhPAJPRravXhi+ylsnMbHgggrDO/3
pUD844qXO4kli38/czzVFMYUmlOyJXNnf/pHPqwt/SAK/9CNgz9YyXgh/OTap6DEhF7s+Ua2vMZO
uGUzAlsukAvrL3EgEZ+a4jvP1BBbEbSBtHv4fF+20+Z72ty+IUq5foWkDp36s4luZlobfO0gwNHn
rsc08L3dxGHO4OaWW4Huvt11auHGAXNEJU/RjWOeQZqszfiy6v7iiWLdNsk7KDUq4lBDb/AHUz0y
TUfP4mnITdmyUhwPi8T5+lWEf7oklizKNxsTw6jf+IofWha/g2DDgZsrEYd7Ob+hWXp/p/vJBC6f
szJvHVMFPB7s2H6TWAAtWBf8OOdebNwnlVXcIqw8XzS9SvEMc+/LYfnTcz9VJgbimRvWIY4aSZ0D
IYUVEyVTZtszJUdIp49zF7oyKTKv6tkgZ4DNeKyiJkIw9ykfhPf1FUU8Ln8augEyvW51M596ER/H
WABYnO7MDtT3n9Zf8gcEWUTzxyYC3MHRQDh4QaYccPTG5RK9WxKppFrAOTnZxizPhh4K0eSSFe6v
rzSa3qpmPqjAEBHMu5kJWi1GNA+5/bMtdTeVFHhakhD/Vh0DduOT+HTriPV9zCVCj6W69WIiZA3b
vX9l278Zgn66vK1EEM55fi171yJcVXqH4pW3poFVmmjJpB7LI/K1sp6xPN5NF8KKL/pkIayBB+6G
N++lrTnmhj1F2ed2DtkMn/eNquw3ZW3KRpsl0C+MyXttJjGzlb0GxQZwSgbntC7XKZWrmJX/U4XX
QtiPXz4AwNuGBjJ6Uqg8vWTjKQzqRoc1Fpie6ZPEX12BJ1qqXP8Ua9N9v8hiDJpD4OfrLuvvLvR9
8r0bLwguEvyy9jEIkIZcMZuMjk1X+ZfS+4H7LOO/NgsQCnkmss49QvQuNmO9oCl7GgvzfIDGuAUz
9R3ew5jHwvzYPYEmipjRKRKe99pebKOx3D7G58W/vKbDZ0ESr0E9I+Hnnd1DlXUPC9KAfwQ68kGm
cc5a58zRr2KSThbHgZOxe/r6wMx/ef7FxeZGU7ovHWqeaV+UQ1rO9lRpwvYCThb0Gulszne85pX8
gHqlVGpU1Kp+iPCsZaXhsTeA6HpVWBPa+/yrSYBv2Ie8lgzW8E1UysB93KUv89OXGx+eGguVfGIM
04VfIs03X3f/h5hjUMZFhjH6ZEu5Z1SDqp6ngvE8QtMlyJ5y8/VwtYudqzLpqNCV7D38jBEeRcRW
VLq2+ilhWedpm8l3lmouTrMD+wSGiKrdfDG51t9xGQnYzna2dExXfW4K2ydlp7iSC0z+BSVpc0rr
EVzQLGJPgFGArc0gQZQaVqtlUs2n/I3BFGFFfWuanHSzqoOwKMWkWgTUyAmwe84qz2PJ+yco5WhZ
KUT3jDtULvtWrzsFEWmk3Y22mQYz5cARqSSlesgy0Y3diH7Xr66yPlVHMzNB+FS/1fiyCOGT5Fds
EbGsPQ/v5pqIX61PoPUprW6im//9gy1r6Zg3PkbEsEzwKMEZJ3cacZnvYa3/6l4PkBEXbeOy3Krc
bwg+Qi+12lEJiibugQG8lj2rWxevkBZy5xcjxsZ2E0v2pYI6GFSy8+Rts8v8br6jF0ATsD+TKUrc
dcsvpERz+89EN/A5YwVqYGCawbMPjwnjg766YOTWoWcC0iZ06TVEGCsxL0iwrTqZXwDM0TehnAAq
k9HDrMdvUHwhYSILNxWmyP7S1KzHYHs0wLTA+IbBrJIBJwWZ0i/QqY3znauqP2ucSDljD8RlmvTZ
8sJLobgu6N6TPGZT729+xh1Z/ErFg7DT8RU6hiwHxuUeDE5PsBn3xL8c7QUqkOkjtbbatsi0UeY6
PaiRT4UZprwV2ITQ1Qt5FhAYBzi9F8zXDN8Am8I1YWO3Wdcp1w5XdNaR34Q2whlRw/IbX+eCHal3
8SZWWSUjWrWC+rJqqB7kyGpamf+c4ImHdQIH9u3z3QjGxaGGd9pq8eaE+RK7Jrq8qWK64GL/heKT
eCpZBQvuD4OG8Ufpr7RFsacYjaUCtnyR74F+pFJk1tzAaAXmhsqEiNr1JSphnms6Hymxwoapqfxa
RImEsb1F2ccxm0jF4olTdgqNziFJPcGspXLaKyDLLfIEdP374lBNEb1QVptdzH6dXbTs9YSKYaBk
YVZ4e1u7K1WgT7EXPNT8Clx2bYyjCe+adQUyBmqMPveQmcHoweO1P+tQoSRP4madpZVoTPtN0y05
WtrVjkNJQM6EAd9SvLx2t2Dy0SJ+2PfyXEbLkz2ooimSbReQV8coK2ALLVp0ADktfpZ6IJn3mky3
nAVGxwcd5T8hDSYTtOqtHD8XokAjiy6DFUfIj5KJpvAaSW3tCee2Xi+rPO6HWkc4VB0EBZ6ZnxHQ
ZrZEm9FlQIRcO6VSdd7oGI7goMgx6hBlQpl/73ZibUK0nLoWzfqmE1h9va2me0YbwDUWoU0QK0NV
lL2W9nDBNwWJIX1Skro834lZ0GiWILTDZ5FYT05NMQBmIt9HM89EOYs1473V9AGd1sS0PgL2s7Zu
3T0bjj3sd8FTHlghFbYadeBAXSmqmmCm+laCNDKgaoShB1yoaFpFc/iGUAktUNfvfLNGQmbfj0DU
Dl3RqJErtig2GfrsLoHSXd4zg75So2njQLbonffxziIqFXwVHPinCizYCtdzYxcsmg/OSfA+Kfci
gx0yO6W4HiaZem8JIlsJeeK73HjOfPWq6ptSpsbCzJA64cv7ZwqCEqAWXNxAilAJYuZ1PE2Khejp
3DQ8aYZ6KnpwaLi5PDPXgFHEVn9mQcvSqAzkGRrD06TlZKqgZvRnU2Mxnerfb8ePiST2CLM/gt4I
/ieKx6Gk3QaDKqB+ztoNa+BGz/CajbJIGKnsAzcYdbXcVtcFuGbmHUNtGQi93+gnlLqzUG78A/mi
aoHoLZKtsRWtp7PmyYlErZF+/Lio2QvSWPeej/ij8tyY3pz2/LPyMWB8nJ5ayseCU9UXz5N1iGdY
1Ew3lkCUwxhojxzFOpl/SvHQuYIaBOhOGnDwHPN53iiObUoBJZr5AqKDih9IK58oU6lpaFEKiyrQ
ndU+595ic2o8etRXQ33VwgjupFqIw9fFn5f2MxXzThjY9Yf/OFRgG+Rp/qd3Fw/L1xtt3X9xTNfZ
wTKUhYG4xq+h9F60oiIBG0FWO81LyXg7ZJF9wjZEDySscnZbzfkDInlp7TQRygftISILkpmr9xbp
KAh+O2a16TRo7H5YcfnU5Uo8AutG8R/plbnjidkASVxyz+ltMnPKrxOo3u/yc4422n2AZ5Tsy6F+
ONwNWrlX9LMKgGgH/dVmM7dVSgumOuBO5cdztDo9xYiyi38O5Mga+58dEP9BPC+v11skiVAWm4h/
KSVl6B9fl8M78L7gM6ZPpFv17NwtzvNxEKwxPHKnC2lZ0QtBFYyHsZ2E0RwQGzVvLYfmSX08BKfB
ST7TVFBnbN/HXbQY+hXbdStutrb4Mp1138hEbZXdkUFeIiDfZtgTFuPLzvctRZZpyNCMD9KnN/so
7JpZy7REJ39tW/r3OGO9gFRQVbkLA7JVzRp3jaTZYMZKiFnO6CZCthKKaYuLepNQ+MWWfYAQSnN0
w0hv7lGdbM66Dwm49n4k1Z4Vcwf78r1CQK+yNEtSaY7zunX5gI+s8gj93pqPFmOCMHjfgFRyg6M0
EcgAepBbafUa3imq6D9J+2tWNQ9IYn35cn3cfeQD7Y1L2fs2/osjTxeIW2S45JE9c84iETulsZV9
Tlt5L5OdPn2hron/nOVv94vgcdVXINRC040jG1rcPw70W9HZSon4v4GqFoX662G6ZN/BrY7DOD5x
JW4djvd45WGaOlFmBJR+RX9djiDR4IgXg1rgv81rv6grgvNgZIwC9qbBTmWSjr6g3RJjWMHWpVkJ
FBTxpnYOiyb5YC2fpz0n94WeSXYqNjmGhrQdZV/4xw2bRHmmJ+Q8oCmiVK7zXUENm1hXd+J1ejqk
r2EnLwh9HSo3qD7vcEq28WLue098ZvL27R/wm7vEFQh1i0HDhZr+/uPMvoyi5iKvQkOSXsP6sgcH
OLn3rbSIKIw3x5nBeY7k9NmPVisItO3jOBY3toM2w6ZAD7CFLVBGhuvv/PcWVyuuuKZbsOcLoCPC
OWcmk4skkALoNmKD0iL3F4jtiCabd6cXhz8KMiKfxfGYCGPzeb50xSWj1vCIO6ISumkC5HhjN+16
it7xkR7ONj3FFrkA4z080V5yt2cCkpCjb+SsiLW/2E/6E98lshqTtk6f8c5yMmYghFQql/1G6UHv
h/hB/W4Ooe1wpP4Jiv/kfLH68SpEVAXbPkVNUHEBsHKQSnHt+XqOHNj830WVeArPuAOvTpoG5Rpc
kefbTyyYLdE2zln/3jVHgVIz5G53AhxG5gy+C1g7EKNMZznf4OWgBHKEielb7t1ENceOLlG2lkJs
cje+V71g8JgL4OxhU7BOv9YZlXSWYPTBUzre6mKpxNcXqUtMgOuRhcwf9Szc2SkizaAl9XykrNKp
x87NOovefUN2HHeS/XZ7CIg7kFxByHmsaXjKQ3sGBQ/htjkPlMnYiElzpvWYPnQkoI7YonRnrQ78
uT6hebjMyo0HUxYE8SHJv16aGJhonXURhzTZH/ky8TzNwm9sgfU53NDA6WaPgskR3h6GCquI0xcY
W2bmzjNHFEW6L8vw40iiUGuwjj4raPPqL/jMMdVI78NSZUsCRzhMGIbek6u9LOa56RXwdLR5ICCP
XzmGo45YNV3Ud8bj0Ux5W5rK7AAjZDHKaT7D4ejZWkTiX1OgPqDBjZFcE5BPFcLK6oiWjzYZ4gPh
uiIqi2ezJ7MHp9T32J25MSfbCpMuaTXQFYAfTKg5Zwa1uMykFc5jagjPyRPO6uu1sOuRFLQcbuxa
TnNXxwKPBzEmTf1CPVgimhhcTBoZ4YRqa0s01ePosWaTRkv6f92RY0VzVXoXowtyZ45k01bu41CE
eYrMxhIF49iPWKmPQ3K9uFvB9OJk7pANnahGuzSPS0x6K6+ACg7ERdlwefl4zMwsL15GED3exf9b
DtV4HVj6geY7O7vhZyYISISJpXcc7tF+dj+h924wkAcHqQVzs0RN2TIkQtDV6/Ht9+Jub080mzdx
q6FDEcZqmO7TUCqClWBaH6WKkvcQ3Zjnv6kdra5hdG8T2L4LRMlSPqFs4VSUQY5kY49Mx3qdij8E
luvN3B0GlEgi7YSeUndeCJxnRkZOLDe/q3hp4Xj4PpKkck7mtuwyqxdODr5My0YUZFnlJf4WOLUq
/U03iMrxrU7yOP5OJvYFuN/mZALHrNJORKm/A7M4sjm+o8eh5m7uLq+cE3OV5FkZ7MPf+xRMISE5
EN7l9i9B9aD97/+qgKoky1FTAXkLci/o27dNu7SgNk0QPtQUxXVo75jtpCeOZ01Ehl0+AE7WMt8U
8U4IuT83dONZe+lQnkKjk3XG545i27Alfyr/AlS2wJLfczWI2y6A4qHrHIX2Unb3LOmxGsGKp2er
tZSeGzoGycCmfleX4MfQc1igQt2+HIJMRnwlRP68D7cBK0eOd0hLi2MKpFd9G7FxBfM0r5GtzOMT
s8Z9gM3KirK5I43YfPg0EUthnMavjiTyo6M4M9UQLPn4Zes3NZzc450PEiE8CTON8LV5rt04HaIN
+hxZOpAwbB5q6MrcDHOIL9uco+xAsgMVtmlJL+PPFKncpbEQnCR6jqsBMlDpRz4zfOMNe7X+cddc
jMvHwJ+sJf4Afwb2Egw/onMxxGTPyH3hRYMuClV4XeLRuvrCulWmQTGRhr3j0rH9hEtl6CZbpQi1
DenQjk2QtB3ARnmy/d/Z1QKcc1lV8leoclsbjChHXoZBqP0cX4SH7QENY+hkjoydeEme0UyfLv85
85Y4I/ExXZAiBLO5giY1V7ZHJBz5aAi5LmFtkPVfQ5dFINHMJ6Rq1y/9n4IE2smrvvpfwCtGouGn
qx9ti8K8lIYitFUQfLF6LRu799gf/sFC2gPDNOtMIhBYUrdvunSWc522sZkXApEgovbjYRjkXasg
KIgwQMVtmrimZbpXOYGwl1Vm9oeS2DbLN329AV/pGjdhOSUenyAl8RCw4ruTK5cm18FBc+n152xe
2hS8JR5YpPCvKvLGGdX2MfGXdzx0udY9oOcfn06zjBCRduMhE4L1wNpojntmWUUxnxEuTUgjV6Ei
Xa3VjrHfHzLypjg8i6hGJviMtD3EvBj5upsZJaDTbV9arOyK0ldfoBV4MREKGzWiNvETtAqiitt0
p5Q/yL/wz2OzM89/iZ4PePSVBkppteCow7QonIuiNvNGpSXToPSpsEhv3stcDujYKI2FMa4NdwzM
H2BnspbMLNnP0b3vQqKIi4fr/WhcpL+bm4+fpEBviq3e8IWZ/mVHe+S/DIgtZMpTfILP/intFzZJ
SZbzxOimi/mTBMzMYmeKmgY5xOwBcTXeyr3GdtlhhfP9NprlHNemVu4YMrhPsI0HHNKXs1ksARxr
RPv0+joH1nIPwacBsYXNOKKcZkGVDXhhKN2rmfl9Ekh13ye2UAx2mfK+uhF0Roax/bR/knNIyXtw
4ALrjT6bBi+VBba/vYt5HuykqphlWFcbdamdhRcSUrALZmLMbkc9/Wj2et89h7vas9cSNwjadVC6
JUumcrSRlTno6fV1DZFl21mc+gh6DoPASzEQj0g0mbkVhCF22T6i4JEPTt7SVnw5o+GCcxjTyODd
Ax3G4CzT+WA2OOgRz+ZkXugqErwcMFQc9qs2Y+/DTYvLRLEKdv1isNkRx+xr3haKP+uhwe5WxuUg
JYn+9mjYvzhYiRBz6iG+YcKJuEb/m8Snz/MHo1qRNXYtOG9Op9zAelgkNg2jfb/VHaeAeElufX+x
AbGRbl2ppFU/PKYLCmZZxxXseXmkirBXAj/D0J+/Dws5bIXc3IU9VU96Nep/jYEiJ3BgPyK0Be3F
qTVqDcWC2jZ07gZWoAy5WfVX9mPeGu9+iSLkhNvySUsPdRTscMYNqrrSfmJCO8cFESHjDYp+hDAV
RJPvnv8SfgCPYUtZ0EG/IEJ0UwSImx8WvQp2gGRmLHwciVVlg2ioElqElJDmiYGmmXPxWG7Le3MJ
TlD2qoW23yUdtq8ly0AnRKN3QGT6+SPYuwrs2C1qTd8NKodJjytFaWBEdm30IBojLXWqUDGEQKxc
eps4HrRT0LgqsAPbmmQSKeW8SNsDy/wwI9ZHfSY9BMY3ehtzQQyskCoIDWZfUcZiApS/+q1cHyJw
OrDGFQjnLquEtTn1gJg9sIFN4wbCTPGPc8VE37aIjvvrqU6neYdHkGo8PJOPn1YhfDFGTjw6q9Cr
Kqx0BPz82Ld0lPx5J7HjLuUMbs9PQcsdm5f1PkD1qzBOry6HUfZxkOVXoCk+AOY4Vidj7T1uDDD8
FzExjevS9j5nFzWdT6lmR8MLYvpmITozvoMXomcnJ9hJ5WepwADPuTlGpfBROjsvpgMqUshovISn
t/qyu5UsijqwpH6y8Z3M6WDtpFe3oklTDLfUJh+XO4uKvwC6pqkVGO88CXHhVp0U3ZPrVjslvjdb
rjbENydOJg22m+7fWGWDbaw9VVp2dul+sT8N/EqLq+hj01lhAznWd2B2SEEhR5uJY/NpgqBDuRzH
tEtUDjSoodOkVrJzY42tcEP9rMxLwLlk/mKMyK7MpgJ7NzEyi3l8R1pw0WU2zYruHobjwngWUgMD
cpEKmw9v4l3U5Y6Prl70pg9MNw48aI3mvOx7MueLYUzCYV6fboPygP3ydHmrjt/7RYZhfMAQmK27
8SBK19bCfvNm3dnuins11Mn9dFBsQadCoWdUnEd23E7vuemyc+0iz+EXlEAicN+xyFiXRmW/zVcx
Cg763KFG0LD/TnQSIEMppeeYFR6bpC+TDZavla3SDQZ/U+3LJvNvOyPx60N1NRqsO3TYDl10qaNq
MaYeen/OP3Ptm94A27Qr8NRwWxC1fVOqoOi295Xmy9CoNLaaL5kpwj/7vHVL6uo2BfPB8hpYipxL
agQ57/Eq8wM9Ff6GiBZJUU0snH/l3M8H1y769CLfqxpbtZ85dRgW1QGcHVKW30rhXSx9hHXpN0wg
+VftCLX9Yp4SreWT6eixQoQAA53SFn/t91MENZdT9RLfdaJ/Ov/rRh9tmUY1P3RRhNFjJ1zJaD+d
ok3czbdyaVCUcRjI7lUGa2NugbVPVqY3dhdx0YyGeknGA79lluAVV9VZ3CnKbHNtHe9OqoxAElqO
owCo4RBGWwM45FO5Q41sXkMMCeb6CCpoGM9P1w/UiFgN2UIye7L4CfAL5opOkumJ3SZpFAKNMyE4
9NE3ZZixGUGZ1gnFRKFrj9LzhNiNpd3hcDn7cmHJ6QOOAI5YmZtskorHNls/wWT8UzOYrbwA1DoO
4tN5uyuGXbQhYSYpEAfGk7t9IPkGdwhTjCyrYy0ry0mkeRODRsm+p9XSQ7Fo9K4VWGiGg4/0TVr3
OsFGB8rbzt7ED+gJQc6l8Xb4BoX67CRF9njeZFQurm0BLSl6uqcLFByohce6JOvQP3aLJHMzZwYy
oPJOx6l+g+I7IZfBYNe+AJN9kIvOb+vKf9PT4GFh23xS3B+wK5Q94ee73AahevdhysU1s6x+tzBM
q1A1VR3DDaXVqqGqjmzEv3NzoS5w30FE6BM/GubwPDHDYpfg8L3dYoZvNDw8Q4QhgpCeEHraJjAn
GpT4NuPWLFim/0jpLm7XXV9JCTma9jj1pUbrHdHkxLp47USTLKYTebkE8S0i2CashidzBzoVWSU9
1eTqEVA5p5tWj6cfz/nesJqCNo21Dof0BKlEcXwwWDvqv2sTL6r88peoUxSLC1cgCJI4AG/mVrF4
bSP2HubQgCooakyR/JPRpxwR+DxuUPsxQK7N1Dasy/nUq9WasYLoj2jAJRUrMteGuElhvWCDIKV9
CfaSCUI8FpdAI2EMGdid2w5lD5E3tiZ2D8O5OM/iAVunCrfOJzHmiD7siWuux9KgA74ylorefboC
dx+udCcwbqANDVGY+x+uXeODv/fLy6C/fH9D3gschkl86Lwo0A0aNEq2mfsp75acHTYBe605NJ78
HpT0OBCm95eFLMJN/9CthJ3E8iU1WKDenLlNftaOowtLXCWWaR/ClO7vldYprp2IiYPampG8UifJ
vPtbuWX63PHVjY6rCSqif/Kt5zhit34XANVG7s5dBpz9LPBGS+z0RscuYZzrTTzF/qsGSYs/ZuDo
9IaFV/jvQtglyXQAWm8kZMFguE0vDfGIGSVgZesf79bViv1b2RWDkGa6mZSRVO4p6N7+Qh4oWs2a
LOJm050M8TMVOdLX/95Juy1QwSeCxZDpp1Io/Scz9pboNvtFsIzef8Ami3V7K13chvV+ah+RYp2a
aFHgmuhOq4UCjkzNEKzslneym7hN4KDrpWFHTsd/LO7cMOpz8lfGgmHZPi8CDN0SljrVJQKQsYYj
uDRYIWyFwZ3NlUTEAvR6y4Dv5f83Rw3477wz6R76y36oCi0CA+yO3NPcyBfw7BP8j8GUrsQaxEoR
S83VeTpk19dVVoslFpr9Fj+tsoAYcRirk0Vj7El7bMXf7tV+SV5y9mbIEPzytIc2LFkjqUgMayx/
ft98TdQRXE7PdYqGLRa+Hex1nBOx4uBVT7CM1+tZlrU8lL8K55uxTMJFJgdmj8JkbAiibyOjMJvU
BKyP32fXZlFoTYqEeXrScod6po1EFMj2ctFX3lb2AZd3kbxMQhMHAww781+tWIkdm3HrMTtsx65m
cQK4U6xR1VW+pJDOQhPFj+L4hKcidsoKpn8cQnzHoxqLqFUvSxXSYqWACy0JEZBPjFmoz2kKQTMz
wkbMWT+/TQoinkkkJhFpQAPSFN3nIUEG+BfDRH8RXE/+DehE6s+YKLbyu+nkJnMiK5WoiY2x8Ozr
Kg7QX22EOQUgFFHcqhU7aEmg/kW7R9Sm4Zfrs0wuD3Pl0IU2G7Cv2QeaM4We8/h5Hxg8hlbBj5v9
tu8+3sKxxLMhY+h+ozzDX+lKMqk/MIqPZeuBmJCNEJPRUskxFrb6UnheYXvHiX75+JLH40MPI0Bj
pWl24yebcJ9pt+XGu6zoFe/0bx9+R+Y9KbCZ3rTfIJcxJvCf6ccdQWFzna/r8YIbo2csMSzLfblW
AlLg5e32MNm4x/1ol/u8ZGoeu0EOrdB1OECUF749sddqKVmuP5JwlHnzrFpuOkdu1INvXSPZiH48
JGc+QiFXb7AXCrUFLIIh7ayo8DHSrdfcJgh/VotxfLX5Pa8W4sR84Rcv1dDW0cw/yZkswapxdMnm
+TO022OtnMqA82ImJs0ZR5Xs+PJClTzvtjR0JXE+IZhqievpCxm2xbYEn1LB/CrQrkv1uxwsztYV
n13e865z874b84agJSAc+lS50wBNXbO+yp24j3lswhd66lL0IzlJoP+xlYM/ha2VnhoS2q2DnYgO
HRmc+C8k7N2Z01NM7F7sZrapSZkHmSiRvg/ulH+sIstW3cTe/iSsMwfTPqn5jxQ+sqxs7ctXWwGS
IqPBuwxVUTGs2Yj77rHkd08hsludvbRInNGEtHSQrQpgE5APwUL/pDnTOHyEH7FTbLaoh0sBlKUG
Ywgf67a7ve/REaiMRo5cQJFYboEJLWLsV5O/UctGfo9LxpQPwG3owhhXQ51kZrR7aqSP8M6xRi17
hjaeXS7g4qb01sllYf7jvzVQR/Ll5AjN1gXQTf9hKM2BW2xooWoxqYaSi7J8p6T1vRCOZjnzmZpf
AkEmJjX2XzeuK3CJbn4fj7vFoq9chalre8czIVcKiIAdiMXTpruUbqA+DAY/ll3Zuf6yqsJoACt0
/la4HRRopqh4AIvJHIKyV5hxY2d/U640enZoXlfzRZds2tJ/Pr1qYyWn3TxwvkWz/Jaz/aLZ6yei
h4jlmets+V9Lxpttz0diTKUnNRPGr4vGN0Lq+V23ucfvSHHm07MjhfBOICiDJthhyPcyPCL4Y6bt
oTigibw1cvkRQ8T1kExE/A6MoIBWZlYy6OGxHRFZQBcjV5q+dq6SsilSnnXOJ857prPmuAzOyNrR
JuxJW4QApvaBqsit4Ex7PajhvQpdYkNevzI9zdZxiD2t8ItjqGXor3BG8POVoWxLYkr4L2dRP88I
wAmgsMk46RLfvS56hmCHEQOCAAP6JKBy67vlI/YdJS3puZxpgzSevicmxzS0aViuNTr+9ag4BFeT
7MPM8+1dfCVCn2WFee+SedttcwnC4QKn2sC4nqVJysVH9aMhnODA+8Jye1iOGMFQPbsUUP36v/st
AhgEFeu/H9lqyhYrJiY6cNEulsXtK8P+IF0tHGofnV/0BkinnUD+nXeXk5T8qnf/HhBHrhaAIBPV
hvTnCAxYj6ELoA8e9tW9fHS1DbYPKXtR9qODvjWnsmMo7gcf0E9Upm4hc4tEDt+ss3SxNzjrw4+W
mwZAoUviHxLAjlhRkmnFYp3kkojKu9fdTVIf7rSMq/R6JHTrNh3I/J++KcLzAuSM43eOK+abS4Ue
jTFVZT0eCT0ebwD2vDir+CZ7rCzv0ziTS4A7OOsHmQt9J4XxnkWkbVWzeBkBMUjJJXfLnR5bsPIv
K8o/vXwof+dR0GtPbov8d4EtHdiFvqHHbPSefh96u7vM6ArqKZJSUHSvq6i1U1KLHhq9qoGGWiNy
8F5SeyD5gkDGRFJYLFKX8+q4xf49qhfnMNNU2+N5aHghy9/R0+8jjmt1kZojFNZdR9TTIOalEIQs
yYpSLdYPGEqdqwbFwEhYlXBF+imC1H9c549VfUk0C8nDyXVgoHcZ8cFJdEyh/iArHpJIbIyRAUna
jyy3TSlm3o5xWVKL4zCRnJCFa3iyozYiSa2vE1HStWWXDDw5q905GT+6/FiyZutIpMU63rEDfmkW
Cxa3TvTp32gkFBFBvexmbnXteTlOjK58af0p9VS8WXnA4C1bhCIlRj2/SCoqvHJCtqqWxrTTxpQM
g7b2VN+tOfO5culI40512Gb5FYfXqOkpDgszm3rbjQXQ9n7ORiV2yGZoR7+fLaVY4Qm13w0aTjIu
YAbblakxdnKFIWREREKGPqzVTfWs2aN/HgNFX67Y6Vr2LyOYqG0qd4VBBirZuGOTLle/YMuOrnC+
VmeGncJ3UYLf0d/7Z+EKnZIns24IY/Eox1fYSSCpOv+h+qrDEdLNg+p8gCzVfvcG5Sxu/PrJ7i56
kZl5fOy20UCZgwZEM2xNrWcAVtHmVhLqhDK+oSXsZE5mGExWHNWCCXyVF10OqjzbdhKEdm3S32QV
nmxVEyjsxziuHTNvzRX5APMxTJd/KGsS2xGH99x3EVRNU2LAQ8ah/K6SibwD6goivGpxUP+esozC
9IWF+VNjJh+KhGqg8IvkxeAKbsSEr8pESw+GEzZkaH68FQVww9dTCVGUfhRPEOr2s7RRqy8FHTR6
i5K+inX2xQzXxjs/jpx98X7nz9aTqVFbdW2TAVC7aTfRufsEE6BwU+E93Sxj8INtPgKgyYnCd9IK
ZLKAnYx9+K7cDRz9vQWqIrT+Bcjw49b8znF8atHTi/NUtp1BxpIrQomax8m8in96X2Jm3cpFj0cB
zEKyfe7J8RqTrkfsbYdzbL833Yj2gt74FVNpJnYoZrBUfFmLszOTog/C1WL1dYuxEJFrF3iIjhjr
+lqu0lCOSaoR/HNN1pMSPvHKWMcZaB9J+SBQBE4FSGXARh2sKLVJCSeiACRIJOW6KbXWejlvvNgP
S7OdplxbUmWlpkMwog+EWkRq4SUfQ7DbYMT6sVHwli3QUqfocNsXwd6124Sr9YAOfWm/z8g6DmEK
4UaxaxDraVhg7s6KY3j2EAk26HqSc34sBiwng8oIoI220k+JAD0/+GlonkYAan+ji7QT0JLyKvix
7tWtZPdEXbtqLJWXDDM+nHAAjotE4Z0KfLWpwE3PYoY/H26wNqKz3USo+w88qf0PSiVXWAA+ECEV
3W/quMtyFdiRmQfNTycDzfHP+OQr4Ro52baxMRNLaA/GPMXKvH7UneOBYFcoQFcFdmm0ibgpOsJF
EBJuuRglmUAc2Prs3EjScYz6I3TNA6RQj2wFsdj74QYf1CmlGiPC+E6wGKRRTLjp8aaiQaKYs4yb
6u/QcNBXkx/0nHm0xIMoRqSrMr6v1i3i/9u3fssPLVkTtNYUbazGOJ38A9GmZckYrVI4Z+gLCwJH
J7O1/myX3vkTW+i1GW2UTmzThk07Mrb4tdiK0k42tiaq58HGTwVW5ImhG1U2lV3iioyC5lh3HDR0
iy3oLQQZcj/FzlpxJlsgRwHSCTYyvbqkoQnIrRim2AyJAe5mBirTAdyDQl/plgyuMtch5EbWePD6
cyjKQS3VbBTqIZ6A0GgwpcS0o2xbLvHxQ+pEOOSu3eNSHjwVwdZbC7+1VWqUw4rwPGq2I24l5UOs
4A2vKrWdCgG3fxQ8AkNyXxW/DNRbkFBaiDF1BXZKW/SOp5tVZsFjzbRvmeQj4JHSn4pNPU0IPIrP
BbxtrXcQdHbiDCKuj9KPKms9roR8BHBco3vB6OvsnaAPc8LJrQTqJfO9FERx/V/8Vm/Oyxw6zL7W
IMBbq0a9Dl5a7pS5XkbzVq0AU/sg/pq2ou0v8zhM/l/J7Gi8aH3O02fWnZ4FA9/k3Q0kFjZIue6j
2UK5pG7xv9xXPyBlvJ+OLe0sVHMIzCIvDiy7MDxUszE5gBFF9zlKr1xdiwnB5EtxavTnT6THxEEU
zmfZb2oBZ6fs7u74PpCQMXoB2BEh1NpBFvQ/P0youHPTKEySC04eQwOxnvSKWhcRrv9950Un4ZvV
KUToyUHltFyrdUDjbfxfkOpSHZmwW9yXMcSr1dadfZc0PNnFWy7zpenAq2c1aUfd3JeYYtUOfvWf
eMMnVM3YljtTPC4YDJet5YhDowjhnEu7YAwTeTx2lCQJxYFWKYe66Csa3975LwIqBxGG62wMdZYw
vbIltNnvBIdvqJRZMisDHWoFYsFExWMfdk+XM3cdkWMUwIS8EpTBO9LYGQ4BNZKR9a8OdknA4oBh
pLdUkKdxJkSQbxc4EDsQZXhrkMkzaKN0yV1ZVPwKrxpKm7gMz4sY37F06QnJjuGr00LXKO92dPMh
j69cEIqEI21ZpDQ8uv5NbjPa6O2VFiw+AiKocmw+cTSf7VzUtUkDAK7uoYYPCiMMeQyG2WAozAkh
dm4T3NHwB+kugZZ7l83uZt6cuWlMfIA1uf8+tHGTXZM5aAjvklX1sz0qKVhLkUpC+OktUGi3swbZ
uUV1ZnLrY53AByYaLXQmgev943qwvnwKLodeBxH3hT8JI+WskdHy9yvlM2n6GcwAlmeITKEGEo/a
253ZJa+Z+xGBYR9xEmtX2C3fpcjV83CiUrMOuZWdZKsRudeDgkj4NCSlO4ZT8KXqrtmav3wUVUGo
wnKZWbxISxE+u2Q/R4gGvkxgJP3Y3fnRHChXqSgh/E30vuUEp2HeDJKxtFwLtwrxSyUaA98GeO0U
ib4zBKY4RpJGIiyAzwRRRBFLt2DFHFBqe3WMiK+XqVRTsu1NFymHRp+Je1f4xqNBEl2dLdw4xvHM
T9sZBQrnMTLfC4mjclmFcaNvfaUYQRuruAZVkVrvcK2Kr9k8WMwR5/dvAuPNRWCvp05QHOwq9fKl
TgqNL1bKh46T8XvWBad83OmCXg5pHeqRzZDYt6eevU2u31qUFmejRMPa8f20S/IbCSJcrQexDTWI
kwHrllsgwtNMVPcmVBINY3eXhcc2FpSB1Iw8sJbvgDcxn52W/fruHRQKriNA/HECYoP4lSYW7alp
hfqakvjXy32DjP9Ihpn4/ecjFPVZiX2f9X56jpUy+FJEtQuLUM62giACWs0hQZIEYyLVUvyfWEbO
jQSl77Pv1gcY4ByXzUM8snNmejyU/iJAubQS4+nJlpSeQf+JtmY2pIKzNQJIXlOIvHMgMWNhTAAM
SNVSUXVJKRHqdX5WFTnBR0gr9HYboT2M+m/zy90hMRL2FnJI7YG7bGaoR59dTKxzNua472LWN5RG
9wky5OCAzcEQ4fEBGEYmO23yW0Z+c0swZpIUXQPqQTRiq3gTR3HY7XL6ee1gVwI2/yYB9GrdQtos
W16kbeQiQSt90jx8IFEHZZ/nuI8+Rw1CHrO3eoU7UwdhcY0jYjUhblDFa5nSdPIYiX+HU2et/fZy
+75FjAa9rWaFgMRstPV1z7EOhqZT7qQ2P95kIV/DJBcthLz0Qj/pdrUsnRqLQiXTKnDq+ppuWHAd
URQ1Z3GWBHVQ7Ufh8zvBeaD/sZTrWGJQdYxWfj8ZBUdSFHbMwI9H3a8/l75pIH9OccqthRf209C7
a9+Ermm2qZ2+96MMXcfv6IxcDJo4kKKFF8I65tAdQlg9XC40zJMp7oQxH6JhIK0/PhEHWlCCgUYw
Ugq9t+/tDkB3qdT+TJmSPm0E0wNBdhxRAcBt+cAWJt8U/mNTI1GqwWSEg+vv8sWuf3lTf5jfkUCy
x4itA12X/gpibRHcjB5d08wWCtq6Q9MLNdMvXLcEE4JFz/bgZQFjQGzh9dfZ+sy1AGJV2CO6gqSq
uWI//mNvQuQOZv/cW5Nohpml5WsJt4BHiJjYhOccGj5miWEojVhIKYiUl4uuTlLPMUn3Z4Hbo7cw
EmBgbItdxe6zI180N+Z4IZmS4u3zUL/lDShs4BCmxDATBEdXIpZe0DBR79ka4y7hMa/M14VzJkwD
ZmlPjG++PpkgnS6+H2Xp+1aGxt7v+NuSG1eIyzT54XuB6R/OjEIwvtMht8LlKtEvFeFjTmu0okhy
47g40O/dDVUiNUMAYx5wNMOpTKoRe595F5QblqA8s4Qa+hVWnk2/osOmcBcdPmkSEfZWiSyYz8+T
Bmx8BoPFGyCo9MhWnhQSHVlFNHK076mihnK2XdwnC3CkEhBRxRZOxYc+xnYhqOZk2nRsV5Ur/CXr
IcthRoryijLuo1yPkEHiTvVNHU8UkM12Kurx7Cp8p1YByvERleW9l5K5bADjtyLN+Xso6LhevfGu
0AvcxFdu74AIsVloJOMdrXa8pWYUvUQ4yd1DLG59g0zpEKjqpOo4tHiKA1jv7RakmtE41t3StuN5
vF3LjehCl2PgwOPyqTIxgjcCUYQywBqO9vZE8N//Lw6GTD1oqVZf0om5MLOiE90T4xt6FcG0HKd4
D3uUzcT71hk/c61T77ts94n1rCA+eFbvye7wombzr1pgOHpIr25x+wx8jmseoaW3sOZPRy3NK/0Z
o5WcIP4zHec4IvRAxKoRzSdE/IxOJRJ7jDE6mlMXxChOJt/NGPqtyhPlhr0g7eqITwzDy7g9LaRX
xaa0gqS8AzupBoQ017PErYlpjInFW6zmoxFiqyz24GPiwQOD6kWhJGNzCiCmuM8nLyBrFK1aw2eq
MKl02btvDCgzvgDLA23gMvKAEAG09zqMxl+SiQ88FwCK8SAamxbfLHC33ORRziAQHxCTrxvilgke
CCVqdCBIsf4BDSSXbF3bliYGRg8K9ZybsIAwLjS5OLmxzNUpfbdYn9519d8/UZ2f+ZMeDyW9D+R0
ZVqIC2F2VJ0WT2XLp/UFnIjcg8T1dTmSll+aYA7DrBsz9BrglI2pr6seALcnAVfS4kHGKT9JWj5N
+QoGqayBlSL0vbL4t7ujeijLK2UhqmRYl0V0k6FbddGMBSAYnbah7egCZ1I3/e/ExboVUdSHGejk
iAtAJYS7Vey5HCuUR5ysTgRhRTebbVE5k1iJ2PTxLTQfqK+csUG8KdqcAFfqVoYw3+A95VH+LyV/
26Esi0YZ7U+BImB+vRvLW4dBbOwo9X3kc/OgAkkpI6LGtDuL4dk9lsYRUfTe0lwuM+vsQLIJvoIs
ZMiKFl91w1d9hOijjiPhR6kmPsq+T9/bKY9CNkuTNIzrLrG/L/nDi7oR0fva+rdOZtf470S8J8Ta
MreRc7txbkTCPH9yRK8EcP6a5b1DSe7QkGG4zQ2RbqqKJO9vQGTyY/iokJq8jGSD08gi1cGDDO5P
3oPsEGJ1WWePxk8LtEqfTXnh3MlhuubR+Tz3aGJuSCRV4b2rbou58qsOdaGRN/rfl2kVHZPqypnX
nsczIeFtYjMPoqsBWLzDijBzd2pMAYViBC1ma285bmLWvX1rfqtwpaah5w84n19+7dNwuyldvYaS
FZe2jHqMwpTEJwn/WxrkXwaYvlB701q9ahaoG50uvgXva8ayFXg05B0ffmRrrYxArqAf3bzucmIN
dVOLUXkU+LnDVySMo407R+NrmQWwQ8dQcEVtWnuYaGpKBIUoWRSZ4fZRBSb6Rhkl0OWSQPDloksG
s9WnnfnBQ8r/ZRca5cSw7XgjdEhdIVkFLTVjj0nzdFLquLLQGUo55CrMbZFTF/MgV2M6U3fKIyXS
bEaZR+D5R+X3YhhpLXX9Jv+qzonvJZqMnOGIEVxYaT5vQjKvz2JKepNVgBAQpZSTahcEVpg1H1OL
G1YDlhe229dF7E00e4E7zIxBiD7jF10UUn/qEPLfhn/CAl3yFU+K2c/L93iXFDHlg0oN/78Dxyw8
EAESCP9BEdJ24+h4SY0RhWRmx9IxWrA/i4+oLxJb8HjDvalyUrzt4hjs5fwHbmjsYvQv25/kTtA9
K2TCN/UzfVlR/yOJ8jro3/jwU6b3KewlHWjEgyXEY1qzYi4VQ0ISzQwMwm0YTb5nNA2K3Rxf12I9
WQu+yvCab/oZijnhEUqs8J9c9btyrNGLirubUDc3yk1C9V+pb5r1g6HVyrLjpBVksRgctEeViRdf
RQxmOIrw5hsi/X/L6bS/o0OReSrAVSVJMnpXjH38hyEf0ALMvRo95dvMFGOIQJCNq1Q0pD4nam7S
kKOrGEwBMtRR/1zK5O7tfDwPF/kdcwvqu2B7vFii1h8rON8JzYRBgCtGSwrlGJ46Evom6+8saSJJ
jLL7t5td1WeFmnyGEWFBUhwhGyywtri3fdpJ1PLb00lh51T5jXKHdfBOH+e/LGbI8WTvnB58kBCk
eauZuB6KlVQl5CgFR769g5c9u8WEqjj03JWMKcvP+t+1SELe5pqrUxbuRE69lSrXnqZ8jb/wEooA
+vMMFHYMa51i3ceA8wed4uR7gMsLwfHA8GmLK8gVv3FJeOmsRS3wGoLQXqYy85yqBz8Tqz57SViv
/bZHHtg8nXZjSSIuU2MSzKF3SMRrsDxX0niyJ1in5qpx06QKw5nJa4sa1TxF2zaGxs1AJ1xDpItd
5e8so9NiQasNtISe2fvbMqOb18i46gXXeAJ+4s+LuEEzrCzQkVB16pVV4cZyhw+MHOJ+yUFEZTH0
4J+v6UDGwy7pTdkBMiqKOqBUkjSvoWZXVHKWc0ooUhz0R+yZMWQ3zhePxLjWQzXVrwtB8WMijCcO
zIfw0M68ngOKmnkzWRUfxCw1kpOhDc9KjI9OVEHijyYWHo2s6PMHFEkst6RhTvwukfKqxSTZLgV7
dOJsTyaFgV8KcKYNi2fti/yQv9SZq7IrKhAcValnAP/tEfC0D1Hm2Tfon7kOg91sYdD9HpR7gqal
lAnC8VDjRcxkhMOq3aBI4r607uHk+jWaNgUrP9d26TIbHhR1sAHqFWvuBayeRJ5edgGGsXkNugH8
0QfF4uD2eIoeC/Mr39J+UJxxtmDe//6aTTNOEYOlxNVmEPCs0ZJu8aIEhtbVXIOCVxFKfmWeJSAI
rLUD/gZHKbarQThN1qMX3C2z9r5UqcUKo/mI+ticWjtF3OrfkWQ7ke+dFQZsxINIWBW0Iee3k4A/
uXkcmRBtlB6NQo/3aIq/+HTEZE5E2C7vWSfQU2d/Xhi+18SlYkoSslDkJWjmiSyHW47ScQ2dywzN
OKzNf+8nygvgJP03HNSfS/DKc6ghqPmAFpDXLE5ZunjAR0EzSnAGpYChgVHKlwzrzD4MAGKQvW7U
uz2emLNf+dIsdEatXVjYxsKud3iHIHJTMBzvjYMI8YbVmyW5iTpr4HiJ7rKbsR97no2Mpz3Pbfef
YdfnwsYOx2L/Ai1A5ucpoB7H9D5Vvo6Dfm/b2Zq20exBOkCQvV0N/DFgJ814Cr7HyuMbks/XUyEP
1MUF+0YeURWs5fJuDhQNCeRVNQVqCzJQGc9SVOzRTwYZjzRqzQUVMcb4/YdZCEbrAAsWOnnAP7ye
zfG++4KfAx2liu+CGx+Tu6n6G76Ymw9h7LHcwQqBGDPSrq+jrjWwxZk0sRtnYfw7Vka8yRS2h+PP
YOgXJ83vH+lzS5sswiSW+1YKqgIalOr9rWoFSWstvNAmAgHQSscWNS/J07uegQNUtH43xXNHBjdj
UjNYNNHEqcTQl+SJDsn6LJpf+RbIdcXdUBS9fVyNMs1QQ06EmHkpa4umJActrRp8ypLMZQNMGbjM
jcZ4GlAiIJJZkD1GX7nv3e8AuuTATAfvsa/GLz+rl9b00Sc1C3tYqBBJJM2pN/dCTP21ueyNkdlS
AwMA8Rh0+bZMfEX43wTjmxbqnWcx02M/l4WHSSOL2dlHxgNiNptNFmc+kQXucCgEI7KcNHNeAd87
ZSNG+MVWHOKfLZl0IaHuqVTg6edcPZe1vLCuQyI0HHnIwUxupyhU9yeP4kRRhi/bvj9fqL0Hjxz9
jQt525eYbl7Zkgoiz/6WSRojV/G8o8A9i++Jd6xLeBEMRusKYELCZmGhH7ifynzmPuWBGeq166rx
NbqkJevtcnrc/xjc+kkJd7fD6cGz5wDbh1fWlq0ED7KOqVOJHR7C5/dXbX+88u/54Q7v3Q4kwCh/
GymheJToeEibDIhrQ/BeTJJcHGog9Nj0wGSvI5Dx/5CRQS8LlqS4U6RBfAKkkS+QF89SiR/vrxL9
KpjEB8vzRIjjLDorgoB4/tn8mI4YwcLXum4CeyOjd5Q5UD2VcslgP1EWb4DfqfoStKbPMLK2NjJs
rnfw7kBIPtfo+136VFYZvlKOfDirugiVGZlk97wxR1xzcxVJtJVLCqJZSzrpZWYZc27egAPAJAoQ
oZJdDyDnNsc2XroH1jU+mTLEfiOS7z9Spo1clKHh6oRI36GTDuwD2hOhJNP7Df0eBAcAgvbTeWG2
IHTe5Rq+mMqpLg3AaZv0rsFaMm9VL7YEqNCWfNXFQSC5FZ4/SF7IrGwh0lMLWBs/f+wiT02RV+dM
pSUrpfOIqlA/t5A+uNZB+jCfV/XEB25RxLuyKbLJGj/D2F84dNIQBWMMfFnZpY1UNoF/EzNQM7Yx
qxADB6p3ZR0DcNB2iG8/6F3MbIQ3K9FBDtYZnrzNwdbgHPgL0KzVt1RpBz2j504iGcktm+yvwmb4
38RE8urlvCGpbkNpY5h4COihGG4B1HH4nBjHtdfydyFMu6drDtwmYUgHMj+dDOL6fw2W36DmZ7og
79gHEKkMyUB3tc8Qa71owrqE7w9bZpjqoffXoDkAWLeh3YIdrL0FDTfXh41jhd2xDFc0U0Vc+E9I
FdyyelDclkYiTWltFsUMPgHviPh9Zn6sjwmwFtYXGMGJFzGfOApkhIGHcU2bvIzE6lIW+vz3s6z/
yskF7p9v5Pxzb7cWFL642Yys7rA7iNXOheASAotlfbhidLBTK9Bm9PFpx9n9oLnwfDY4ccfLXogy
LKUfz3P92/xaK287U/Jn6F6xBMJjJDZnLcDQADTMWyduferxumz3YwuKJqiJRQhVkke6yKkB2tcU
EzwFoMz/UjPIIIfKMKx4CBN26THV5xeMQed5eH3xgCNgkHOTNkxWdJPb37ua2r7+st1IhJ9TBrh3
p/FaCTLKKjmp2xjA9xhZkcMpm9SkOfteHg3U8a8th0zoiXzri1682OLg1iHVXoFh3s/9vbkQpzj3
gLRgWB6vGd/ojg7IBnp0pezSY8N7WesBQeu3zr8qxek91/Hgsybnbxg0xKTom+FQgMoD8gIpns7V
nVIAZJ5hTqvMywJGO4atyPr8BLIL2yrSo0VxjWM/cKjKum6TKBMnkIiAhNuAucW7LVo5RH1sLFl1
hSA+BxhHdR9uDZ/ib64h4ZB+exeRykCP/7zT2eIU/St7o2yfO3Ul3JFkRkGPdObx501kRIpcwkMU
PNxB370ms3ccdgztRugZkfQqFwWeG+/c4zOCQRa3N3VQ6A5DVsIngJGRNipIXRQbk2SaHm0YxaRw
WgtrAsdypNc1+omi+iJSe1Zf2XN63AmX/s5EIJxXLdjQH+VMZ2gfkkVfCGAbZX1jN6umyLeUQ2an
xdFEnFu67+wWedw4ic+x3/hUO6APCq0TpFqEd+BZSg0mwM6g4fHsWNCdlfjVezhTOyh9vYxe6k5W
H7zDnkVi3jwYIuWbXl6xvxTN2KsKupOSTRk53nj0/rEqiaan/1/zKcDttvRDy3OkxmCHIEZpOfNj
tbK7M3pFf18lY5ZAAPyIW1YMY1OarL7beTITbqNN2OQeH4rVqlGnjH8Qbsb1XbGbEXeQdDcknNEA
hcQbVTefXrg8g/cFOa3HgZHr9oyvRUmhcx8Xb7KtBHyQDgaURCqkOyC1k5KNYoHmF407MzX9Away
SFYgjCGyTsq8YcCxID2eVOiedjznX9pixR8QF2ECM6Ve3UyQmxMEJt8l2w3255CXFuUkjU84SB+z
MNsNVwRLKbHvitm5uSzEQ/1NCqISkD3SNhnRw0dgv3+p+J+GJOnhY8Ej4f2eBRauAicZU/quVkl/
n0TrHiWCT38IfxYKgEC2mxg0tw9E2mXOrxT1SIHlna8oGL5wy2qJppVtZb/jZYRzfQVcfOfmWps6
pLVx0hEJr3lnmmSsS+w28jWRTkQ4TLWF/UX837pYu7vSmK7ljzKGpbNGNqBsabo31V36wU6P6Q5R
t31qdYZ2QpgWZ1aRfGYK+xFzTyLMUzouVC99KU5qaExZS4NMfbrylZWnAUNAXP8VjKAU+Mj8LFSN
04VBdDcNCvS5+Q/5xElSBQUWUCC3gL4uoHvQZasSGTl67NDbjLIlSPABO4GZ9+Bu7dqqyNpNuY5o
4wLmcDkbbf85/kowXQqdN2/qdO0D+4YFrBHECHSBqUbi10+XgO33bPRdeP+RHzZzAyuV1JETtARe
40r2Y3YT8keyVWCqF0uvUQXzxJ7JgFommp1uN5B3ic1qjXg/QzgnTzJPIcw35rrn5xmTQJ7jUYcl
IEyZQyFB4SNmSvTl3peoUYygbmVbFmPTBJwngsFuwYjjvWji98rC/NqkWK07MOutdnWuVEFQoZsI
T+tGZL1lGT3Gqq6jxwWk+b9ZyvWc/r2YwX3JFe2HzCc9AdY4kUGuseLC0X7+dHd/E1IBn9EnG8k5
VsqLl7j1FzTkohBgUDg399R9ryTqG6oTeO+QDlOdwj/FljRUg9u1KKlLwv/qvHj1byYUF21TOCgC
n5R0hQQOtLyf6I1gddRFiYJH/qDD01t+s9XIcbwsrsmujytpqdq/O/l7xAqGPD6nhcawF6BYiSo8
f1l5xxG/zLCI10kKnzl/1QCbAj815W0VQpdMZo/VS3A++9J1IpBXTxhyUUXvKolwXXHFzkwECczf
Xj1SpXxGc5pnp4pmoUVazKOykxv+zAuXRdYOlHtE0L3zVvKJ9v25qda97uUbFUe9RoRBV8ej1xr6
yxipJwYFLxWs/Bk6TfNqpQaPWJKulqjZD9HqUshjv0aErOr/i9LMecAGMvpmXoID4ErrZ4L+DeFm
Tq2IyLR6sQddhygBDlH5CB027wIoqlxcQXYCMYT5iRLrKOLff9oxpUPjkUFNRFeE0ZwQ7x0+zngp
lJFxp+YdqNw5IHzr531raIPWjqp8G/fQJGUyrM3Co8eraVIjuz+PGx/hLYaw3dulnHXrDCMjMtnP
ZcppdOhSfZIZykCv6FESo2yH/zS0+nA69ZFxmLw3hbsKBn9zzFP75BY4lKd5ILGv447Ntc4csHEO
JMw6YiJbImsVcxKgSK9xRm83ZI/3etg5IwCFG0Mc5sPA27CbjLpVmoGiVyCcGq0LLXa1QAI81ZiY
ybP0MKTOE8nWfHs7REsK996/KJG7kf+OiEhHAMfog5h8/hK/vZ6wHF+jSOA1zZ9CYVqx0mAPh8/i
E3Eo3BtmQTIqo6VxWdLi/UEVtEI6ww7jpy3b4d3Oix/ZErM6TmczXWMjCqxu2mD/DljTz0xSZVEE
nUJwWYHT3xe8yGv89ORMG6IP5QdHRP8pZ8qme7eUEJ3rX6x+T5RTuVFND9XGUZ5fq8filLguaE+9
IF2hhY8xCJT/UBw2vWlT4LxdNMa8T/UHm8OiB00GGyki9ZXtYtEdUw2EyplNX0qDIXkzoH+epbY5
fSWmUA7p6ZHnuuidgND0HPzpTlgZfWyjfUH9ZKxcBmiph6vP12Pkk9AERLggeIwF9aauLmXN2Lv0
k51WZ+/hKwqpu3n/hVcQs8nDwCrQ538WUR9hIR5WtvyokLhBgRVbiov/Xwj7jygWmuMfh+QTB/aW
mPglB3DuNAVb4BFw+G7UJNnGaX5WCgLwB3QeyLHBBUeJca0TwGAw/hyC0gTlcB6ztje7UU2oCstZ
Lb1E8s59NlC5/q7o98V+iJCNwsKsGtPIyf10wEp5q6+FS14ucAJUHj/TRWBIUwO0a8aPx4JeMDIl
Rh8fXCfyTx7Gx2zB2HaAfhM4+ZzLoaMKg0Z/nPWtEyQGMbQ/Q1fvFCuzblK9jexHdd31ac7Bd0zb
tzlGFfsq5PUZuLFAnyErJdHlGBHNbNpL4vCbxcfFqJ/Mp7sXIJ/aSVwXvbpC3wS76gl8JLHCCw1B
XJgU+uT6nWs4L4gFmIFU6HeN+0r7XVaFSRqk8KxHBJjbj6zYhxpiEHxED/1U/98q5pGmqwvrko0R
PzyV66TCEH1StgqY1W6f8qc6zSyT0pOYf+dcXqC3W8eLZQHurBw0QNpwYx57lX1Gs6tRQitAgZuR
PqEznExtlXDXlvlGOAlaNaEGLLzJvTY/Sy8Tgf5UJ4hBsnb9EhCP9mFN07nSBx1U5T59Dj5tDYqc
N6g+tP8bCQuMsTiDXnCI71EPWWMfxCKXuX02/ywLu/MJlgCLaD6g3k1fkQ4yR/cFOqcrKj7hTDMs
eINheCJJdbl1EkgNAMFBV7Nak7eQhk63n6i4r+gsF4KxRTckPz3aS7IgnXQiHbn080lVIuJbbbeP
iKil4lO3BP/2bpKi77kCrDwu3C0PnAeRFL5aYCpQBe2dLnqwCvtm1r1NFqf5dVwTI3yRjYlIEsqD
im98Ki2ze5JVsPJbl9EMQDlI4cKo+s9Jlfx0zYAeQ8J1TpNIkpIu6E+iK7+Ab8KDzAG+IJwRG76o
l+xg7b7U4EMr/Fw1Jv8iX8M5LGMQKS7m9CgvphV8tY2OE3LDxfyYHzQqTo+f7Jfw0otExJ7kr8sv
rbVt3vwZOJTdw9Y9kZJ+sRjdsxBqMaI8yMaSSiSqC0eF60r2Y8fcSe/9YUXnLcdlV7nmRzAVfG2f
aO7ohBRQWaLYDaCT2RFKj5SOdwAicN9+C8e7hLy/jtPTGcKf2z51brPmMB268iHW7OohTLNWOjXZ
JIqSPCEncS7mpOEijaiElk0Z5BfsrpGGc/gYDUPJUq3oytOKAJESgMCxXfmzebKjjHYR5h9bJUf/
WzR6vCu0WUkjEbXbgclmCIeSwClc4vkriGs/AnIn2Xd//aR6fcMj501adt4iwjkcJIZrcgfwanIK
bK7wA8VGxO8V4MvoBU0apuLEOD0OXBUmTfDULNcMr4sFZkMckYxrfKM6kUumnuEmJA2IUY+Da0TZ
4DZnQQq3ZjOh5Rbb6WTr5H2+zylMQ/sNpgHXVf63SjfycrERVB2MMlxqU+spVFde5s7QUvEB5rQH
7JcW0XmxX+jLZYUuYw+XBgLuwvnoVkweAuIenODj49MkmPrsp1g4I2iGEzTZx4PGyCai77GGurzZ
Gntmro06cJ82KjmglV+JDXyx9PeGbqFXc/Oxe4gw+HiecQvT3hQ6CyS4dQ0S2VM3WAWAO+MRXsvy
KCa3sMZW4sMtc2CvtvuH1AvLMlydLLIOCc9A19rvbo8A76ZfJplfLgHZkvJflvi6Z8EvtziGp9Qi
7v4TDCLiUwphm56eYtFQFVsMiTplPC9OB+GOzBqGY+GeQ0V5OYip7WOIpZU+bSnyCiwkOMnhoqqY
4ea4UcfUNhZR54efuPR/32cizq4i3Dbb1ZXUElgCTdfBgrd9y/MVBm3eTN6Zmqe/9VKIL/x75xLi
Xa9sRUbq+Hs7OutlLNXNOJ3G29rFRJ0Levq1LIKPw4vwm/m5DBoNdiHLpVdT3ZCNLG65h1ilzC8H
wnKtG+7t3XMjlDi36F5wYDMUH7X+IpDRvq2OUgMiPAXmUMsEd0eSKiXw2vMIzoIRUUMP5wZ12Gtq
nrgNeV1hnUzqJ7r5wxl17v8+37VaZArz3rNJBsaVxRJCZ2yGKz/6WgvacJVunzk20PHXRu4hFVbI
agm54B3Gn7jv/ChGSOp96pOCDMb+IpLJM1OVcQcSdABJwxhWaIwsqCop5HeS543XtbgdmZ9w0E99
7qFxfsk3sf+NY2R3fVZOLN9Zo6VG002zxyeiEPaaBVQKSle2Za5XMJAPrJPH149JuFtW4n5zFhO6
2RAxM5oCj76szrYcEL8V9E3Y9jNIcTPJj76n9saynU3v2wNUdN5l5ZsNTu13VDLrIOhroV72Enhr
sjHClT9O7VEUkJ2xkPvzjiaxD10KECY0K4AJmHnoxQZ8IJ4pcjZx4dJsuXaN8fXAxOSJNxge+YQQ
cE9es/rdqIYWl3WQ2RLJ+X0yYEZTcdeYVmZoIZpNOsXReAyhUqOK1Y5+W5DCcXnE4fKAO4wjkfpW
FRp8FSXwz2pFhzK1vqjoF10qDbYITWHIDBPVr9dPkRquMfwpyx9MxbZCHS4pyMBCILI7xklC43Od
wFULSbx363qxDydPJyE8KuuwEHDttkl+VPvVhphMoYzTxQA6IGdxkXqA6dNxOdfSBcPYVkVHGqHu
RHkAYuXY7VxVqIqxbG/Wj5St5Wdt1QfyHzeNuuOL9SbYSAHaMOG3M5vd8F44v8dH5BNOevLfgbqL
ruEKW04yPRSQQFKaUv1fctJYfUlBeyzM0T+CXsVPaXlX9+gy1jt3HX6cA6wuPRYxueH62/hvH+50
KIRKdllrLaK0Gzswpcmatw/+vLr7Pfb53eZewUzzj3tpwKegSR+JZVif4UpayfJHwwdkADmXwo+f
pMtf1PWMDhjNuW0Tqm/McLk7G1M5tJEp+TPQaxPWvtZh61sMzX5Jy6D0NATixN5LJeyDVWV/J+fx
2XzIFBtUoxR8WQeumzU7MS5CWT6FNw/2p5XeipmVs5o4wiqsNZ87xw/xOoDjdAaOmh5gTPFG/BG+
bWRknZshgKOiLpGqqaNkA4rHT9vmXIMlmy/Vc7Vg/GZgHzokjFlkz6whxSinmmYPL3PrRd3ItSxw
QqO+SO0IUt+STRSBZKrgaYrMemtGeZVKnqM0cgUrRqQgzSKcl2H0hf52E1n/cFxtF9/oSOvAYiG0
lb6aqouAi2S7qk7z3lH5sckcVBX/+KD6lXiZMya3JxtH2tTAxmzZWWfIYqs1gsKrtYn7fU1VR06n
X0p0LjkTfn9ym0J9a5ZM6PxdEgVk70gYB/bfqZg9hR2yoPAy+8CvrdtSXGz9Sd6A6+gSQoYsYfKn
GMx8RhfRLs/lrCzKK9AFQnwqj1RTK0tar2Uew+crAvsqTkcNfCBbmgEP1CeBKqVZqPDafftKBxq6
Jn2un8lSjBfDXeJzd+0FFCSxS5oH2sf0fjiwoht+8h7D5IkIxbfGscqtgYe9wZCOJ98CCcJtXY4I
SvdK+qTxddlBSEV99yhnsU0SiqlnF+Z4NZZhKf2HhqFvIo+3MrKGZzeGCU6ZlbROJHrIZRILhhlo
RGCV6nN+zEMr0h15TFLElU0dWVC7NWTqPKTGFIWykFiSxdaB4hubG6Q1lfJXz1NH7kuBneYrJmF/
NPzHv3Sahlj7vNMg7sgcQGN/jNbuyUBIQ80TdOBg9hcpgv+hHEgdiKoaQiQ+PZ3DoNyj5ivJXZS2
eWLYhmxlXymSE28BqYASlyk460XTK/AWd9fHEaNehw4e/L5JJgvR1Vw+p2QqXX+XxkOxouf5aOHw
KOorbTCmo1MyPGzq6vRJY8EJK/ipA/eY5Ji7UVmpknfIIZnV5SxI/IK9BsKjMFRSVbASa+ocJH/N
6RTTyT9BO3fLzK7yLWs9a8fTKflWKQZWyfhKTTpukIknEjNwetuVnSFg33gQ53h+/HmWgx7vtATI
fJcYxnNjrrZ5VcvwSFQYj2TEg29hpDb3AN4Ju9DCK9pOkUFCUol34qdCwMl19vLBkjWMpr7d8W1F
PR+FSOMeRpNGYyVQebIZRijPV5WU1CPFqKWxZkzs8Cc54J/VlKrtRyIHWj1P8+iH+JY9xOwMZh2e
eNEsMNbq5mm+IZirI0g4GdIQ/en5Rq2xZ1NN34ZlaOHC9gPvBm3U4lzWBE46CD7f2Ogz1spIfiAP
mOv3fIOmqn1CZdDROq5qpeKDa2dZX+UzL9+EMwd6xifawDZvHkQIdgZCCYlTzg4ri+z8+73B/P78
MYWLm8XE3rvFaL6G1/sQ8+kd+mnOd7n2Jxn5o5xkWkLbGBSHmVv2efQggAOezwX72ntg9Lqe+P3D
pBBj25BnBX5TaDt0umA1dCfRptGI0CyZsXmEzUJY1k1coKe4HInROxCb7vOAIaclGuhxa5NkbLFw
Lxz+4Zvp0ULPKU8rdJFHeDuM3ougdGIzFMPJBMqrcPoPqLeFbPVMWyGJCsPV75IR4rc78MA7I/5Q
JpSODxnMdOW24o3VlvJWENh3ZBQoSQajwcVpIDaQlLnf/C3azXYKbPew/ur6FFDFIWCvdwONfDlv
CQKnEVz4Y/Quxg4crphiHKj+j1irKWNy00eQR7NXrlu4iBRCGsO+nvsWzVFOgh5E1fAH2zBzmujF
U6yQfo52XSKPfb1lTKhRpeTcjDzUa4P1cpd7im687lUnpdoN+9CjzKYJrKA3dlPPTsEw16HBjJeP
B9Ns2EEMWbfOPahVXrcDZF3xh2RMGshxDBz0qzjASVoyYPH8ihP/7HaGjZpDPVXHQfw7A0OvXry1
YuzZSHe3mNzh83fJmWTqW0N3vSk3Vn0ovKw0K9qznVBVXl8R4/F0WNdWrSlROVeK9aR4GqmZwgpT
0qG80sCFKZEIYhY+MLfqZ9+8U44kwTf/XwAwyqzOsP1Wd+d8sYeV6dbUo/AV3TUs34yAy/fcul5M
KuyWev5AOnRjPXbQJ5YG4RP1Nx0aJD0Y//X0FCpn3ZgyCZ7hW/ri7dCmGb1QiyqprIg2Iq1xQE1D
WVFzPRfQsPxlm1Ia2udQ6yQ/GyyOn6W6KjD5qSnp3+nxzaGcVQLKrIClT7Nmy7AuPeJmkZtWXSZp
RyoA9dzVmHI5Xp6fNwdE6KC+yii52GpiY/v9Lh7K50JLRBNyKOVuG4GYUCBD+FM4nMc2emn3zNHo
po71E3M69YPnYM2vtxJwXLYKAN4EZoSUhI7JiQaLVMZtgJqLBP35K4WvQRjqxivJvXEVSsDqZ5z2
wmmKyoXGv3y/sxr6Vgff5K257mh/f/eBYWQ5PaTwZdne09MyHUF/74QZgtYrSLFosDTTypT+EASZ
KnUD2734xbIKSw6UPcxxnjFt+Y8qViu9n4l9HsSTyA1qpKAyYE4amgoPGC/r6yjTS0hAV7drrYdL
cyd5Fmm6MBZra+BsODLz3M/3FfDudX3n7C05HEbFitifGgIbyruKBHHRgdRMzb7ZGTEZVOYJdIwJ
Psy1GBp65vjn/7s342wQiBtXmqIPO/QLQOd7SMFObxRhjZIe9znk7EvEYhTrz8MWYWDavdmPiXzu
Vd9ThbIU7htLfoh8/EAWTA7FI2CgvkMkbL9vNWf/yw4Q3s5I/Y0SWNGUA1jeQabnG7+NfAgBo3E6
X1wGTuaWqKX0X4y+OV2dkKKb6hF8UcIy5jVNaYExitkB0MWHmq3sKmhUDJfkQqrZwITotrrxYJqM
6herdYxEswcF3h3EDlc0JM9GvLaGeYDewQGTiMqGU0N2c5PPYPSb6dAKQ4HSl42llnYn7LnOnyKt
fBGwKI2Q7WJmJnjguWjzl0xxY7rbty8JzZPa04buieX+KY0PEnqVHCB3yo+cKnfzvXAC/lybDYKm
4gv1POZvFicegkL2KnSwHvzqMWZaeGybuv7DPn7gV+l8eJJviAzaZ/T0VSqXZ8zKNS2iskVH6Dkp
n7eQp6q1G30oTbY8IJj2//i94GPdHQPlH+nRA37ecSPYbcfrguuq5/0VPa13FaB0YU5EU0eNAjG/
8R9m72UkEHsbNKb7Su0ln/jj41z7Y7KjZldYUsgoFcneXFeiH4AWR3YAyyx4np7btvmE7RgoMQsn
eof6bOZJJFhN1l2i9efXvkCVufvGcUeTVABbMghFKCZ333ehh96GktqyjhlBNrmE0abLKvchW5hA
cyHwoXusSa53K4h0Pe9fVvEY7Xu7wF9qMGNh9Mqt5VffYRulToYJXRgoddk0HBPrlaDa2xZv9Xq+
IT6av0x4ga5CG6vYizRNY0ziVZA2wJu+p5Gbv5ygdPyVGqFglmcyfa55Dm9LupveVb+KJ2W7x9yG
she/AdSAyZLk9MVQ5OaD6WOHMlLsQ+Yl7SR1Plad+XxsC4mSx5q4VGwvJKYciHMROB/rDzm0nAWG
YG9VeO656KEJ6sc1W+qMa1luWBN8WrrBTjL35TB6yoCBmaS66N11BZ78pfPB8CwW+pMSOJDBJ/cj
g4NZDsN4DAI4AwGXNBycG/RP4vtqC3jUkUlZCzk8tELaobtemA2YwJL2UGVVwkZ/7ginpB55zHym
QaYKeRDcDh9RSWprk+DBlTFCdxEdJ4R4PPIcHISVvguT1l+ng1mm/MGpXh4q2EpYmNlDz1hNhrEH
0p/oNvBMIc802dU5iVXohGE4iX/CNzj6ovUK+UijwbpBrhhCUTDkWSg1B+tzJTlTsBeLpxcDVEeH
Y0/r1p7djB5Oqi/XsbHFg0O70mdnEBsZ+qmrMvxgHafE2D6AyFdshsikZCWbm2iXK30xLadsuP28
jXdiH9cZpCPcLU3+8F4pFm1cxQGywKf+ZNyKfvfkMBRfjWyV3PMe/HZI7mueGyx9gXZvpgk00HX8
XrZPekP6v7O/M8VACulz9FhCvTzUrvjbZzoeZcrmZQ1RgYrEXqz2RVejUPdkgo0x+dm4RCzYQkc5
KJys+a0QfEovu3p8PMYvb6U61JLu5XIuBwBH5kqsUCXtW/6QYDZLnwyJ5O+jVHknDGFUcoy8JwUt
Cm6f20cyN8BRXKCPvSTcJ+wfxHXdo6XNsbiorJzCY/mBhp+8LTa0KRdzgieHmoaTy4IaIByOxpSF
09bhbB0ZET49CcumhXrYAI6VbG6hB9jV+4dR2+FstALZUBee6w4Hog3uwRMkgsFobTPVdoE9xPpj
dzEOAJI8mC0CIyVS+fjuhYnGThiJAG4viLAplWUz5zabY5poezivd5zaqYETnY1Wf5QaLhsPLnZQ
wCujpLiwMjecZ6qtaHBqxHK+XhsuhQF3w++LiSVwzwN2BDEU2xuMH/gfDvvxZq3oyVx5Ei7WAnal
TY5nh/y+rYXdOOWl+S4pO0+uV2j8l0O62HEgpP7yCiQO29srwjPqPWWUYCv8ghgKI5mwEEPm9STF
ZrJfXhmP54Q4CzIVnbZed55eks2ZsX6qZU3AOAfz9sjV24epq/bn2DJ67n0GmXUHcKLwKmKlMr4t
r9oQnB+9G5qNMDhgjLtqSoeue4K2PydhOEpn3lgTDcy4mYr4KNbx2GxWaine7/hKED+AI/5GRcV3
GrK3/DbgCGxHuhSXj32aoUWDjOb5DAcUqewa5d4ZInaHk0hqiuPehtxG0RS+9bY6LRmyLzekp7o4
QKdfAyMs1++qGAgizCvgVaUVP4pSNYJa1NffQnc5uu0vPy8PXHy8Pfh2CwZeD5YWQ1CL73cGUxnN
CHi+YaeMqtqAcUCYxdZNajoSM1WeRI5BSwdEtk9w84eYFFzF+tzkPm9waWmk1+CP38mJb7RVNFj9
x6rcaFiHk2/OUsBLHkRYPwN95JT0MVet8XhSB1/eii4rGjqNUeivv+NO2u07syA+nASqdavvIfz+
l5RoXUhlTKdyLlr68AwMmFBJezOtHYU/VVrz3713idSSeNsq9F+POFsVbJtKDuuLCf678xbi9Ufs
QZC3FtMjkSK7JM+RYYbgo1+k/PsUwYSqXD9+PowBHmp03DLGW9CIzL/jBm5FUEaHrJ9+BcgM5PYc
Q7VjK4j0kaPH0BSSHokwUOzuGHFzs95Nij4uTfvjyvTU0R36TszGmOcrZ81uqfu3uM0mRC7UtZts
pgDtJPAm5GN+nVVeVhG8UAC5qKD+Qmz6W2E2yfK5qYkgLzdF3pz1FHtiZpme6WVzeXIVAAcqL4XW
dsy2rTqDL8gdcyswtcEeaJoQjjnoONtHm8AkbCO90oTFqs0GXqkkIP+P3J9Md3D7C/i+Nhi8oCOC
54Gog2Bs5EvH3u8l/NRT5++bBNFpZt8tvgCXTm/MRoxMsB4Hli0L8Whsp6k9DTKpvT/X8oIZTpEM
HceQGvKd/B1eF8T13Qg5NXif1gZyXNmgKj55B+k0dbJrdkmTw7qoy+jD9Mpy0uktk/PrXJeFeKjG
6FCQ+zgxja/fZFHMsTIm3QZ360Eyb97hLA5/ZT81+tfMHa5qz9FQopv68C2Yqqw/OHpEHqfEmEBb
jivmh++CWzGUIKc4LDccOCVCJ/WfKr+bzOgJv2XauQgsU+xgFpi8mVvEKeL1FvKArdiYZ+Ter0lG
03VmXs4U9hdEnNwZruOvv0oCPvEWdTEWy3eMetAbuVV/JJ7SqJAXMWlRQa1OiW6nqJWPEHZL+qmt
9t8MLFwlpSoUgi6tUMLZrKJJMKE0/G4LjzdwZi7RHG9MoqJWSXayR2nHEXSnEmy2ui7jU2qfvOCd
tbZwAy0ezTtTScMpDdoBBNMnaI5nq7kUZwttMaNrxaBZA1/Xj5xpb6b13j7EamC/jJnkqDIw6lZx
Qld/frVHEJl61U5/m4OfzVcq/Ck/vPUJfhkTEGBobkShtsqTbO7lkdAOdybvZB11YMphY/IYOz/W
DSVLZLLgc91a+86c8e4hwjW4ITxFbT7I3TTSTOao5SXTQthZlmTRUOCbWyjRo2VTSLmh/m14fBBL
TtQyXjuWJtSTDH4EIZ18APTnwq/bYiBn/kNX4PFK7I8kzpagy8dGGLltSW7SQXG8qOv1yGWhi54U
GVOtzmN3jWkweayjsR9rpWsPgYWUKqfpEGpDecxdJ+Y3krPjQM8hksZvX8OutEFHRJVdZpalh2oe
5/PUe6emBqaMAY8g0awxLlKs5DHMbn0G0PgVvdJPu/qPCY5ilaeBSzkb3r8/tj5NJffdt7VfuTJu
X//lFnYC0sCydu10HSUepZvsXQuBnV00tQmHwjQwsVji4h3PypVKD4oxrh22uopfiQF3cZTO8Lv2
2EXeB+o5wDCkBuCg/85X1F0fNa6/Csb1o6I9k56y9rY0FOP1P+gWWhi2x+Qx7vzGNYj+V/xPq0s5
wx/K3ixM9380rTnsu5j2gN7PUjtEYgC//BHTxmyknJOzVL3ZuWgn+6g8CSn+S2oWUfu2oX0hszmh
vlOcy0HVPwU3QHc3edoDUEiyuw16M8w0+aIVZXCrVdcr6IUSiIER2POn+71iMNn7EuuvI8AAeGpG
dANqDGiXl8213OIouIkFMkvpUkRro7GR5pF8aHtGyP4lXFUz12xkUJ6T/Gacr1VstQPn5qxOIwCR
mrRvJ1Kb9B6ul3j/SY4sD5ouVWvgRC6OePkH+STKGgWstZohH6kGfM7QM3uOY4WyTBo+/Wp7zJnF
8JY3XsR61seMkI7TRWtwTJTOn3vhcncl4HtmztZzRlnL4X/oTEECUiiCtLfTh+1IKsciG6C42pIP
QseB4ZkVv6SsyXBUxGNdczpRd3JgdShe1tiKKg/2+fUOOfE2j8KQ0kxKqcOrOmSO1U0VWiR27gT0
LBmwyoGxzLnjdaBba97eaGCOc15+W2Wt53tpVKfKWhhIiZkwPhuh3JkSPQGXeKMjnqZ5Eqaz3FI8
QwR6D8hk/XZY8BVGcsaIqYWfctl8vlBNYv8N/VYBXgneCWoooeHmpRvlCiFjaAzejVtV5zXIb0to
7f5MrsGY02Ozor07t9n2gnvG1uxdD0FRnA7/8MDoxUskhQ7NqW8QhaFAtyT4pHKwE7lb+MoNZgZ9
lXvba55rDrNtlpDf6HUVxYQA6DhuyGZzMHwClgbGOJBEfCACVN4iZacPPh5FJip9aJ+Yy9WY068K
Azqd7LApIZoQRaKFiYf6BH849ZF0Ah3BPJgNK6/64lrbH9lQ8fJyBca0+pIDKuMB0T0lv33gVvHu
/43mU0xO/98uNwf6hhW29uqxa0OWxoSMJkof60e9WCwDgSekexy+fZu6xfhMDXTKqXqu/WFKTS6C
bGIxZSAeexYo6qH8drZrRwAlFBhtlr2vjABOeygwYgA0u5/llrfvRYC/q1Kp6EsYPZuBluPyzBKd
qjx3kOgmaJDg45mVsLKsnxPacbh1dSINDiy/z/tk+Y1mKtgzIRIAy3FRsxWKH3ngBU7Sls2LLTDg
ijgPMsyYDmC1Y7xY+bWyFT8ph2JDZQvfzJ7sTjk1ZSSFAleI/8w/A/YyFCtTVB/2r7sER1PmBwjZ
bszx06M/ZQbA2sd2jmTomKvQy1SfEShPaTUUjRGDc1ognZRYfGLelMyb3dbi051VXy/VVkbcaQ7t
mh9BDYue/5YBCjhJWW/8r6ngwg6fgf4sBtJ+53hfteuODvnwq7IzAodLmDC6gjbBWMfYRaDLKwc0
TDzwPVRoFlpq1prEJ/k2Hj1GomDfCwppt4iXS0AYegNiHQQADmmECr/jWJ1Bx2uYyIFE6JqXCVz6
rOP/b2aemf4AU8aTWeIWkebED+J67/OsMWiXa0zGOCbacZg1/ajDDHIANXDDqOZxXSFsCeheCDWE
VJJZiusyhSZ7+CenkZ8M/oM1uKf1SKX+jVMK/qdI7+nU03e0r01qBWOJMzWmM4EKzzS1usE5lolX
ZcL+nW7sADeEtI2iEOe4nwUt/tlyAJCe6npBIDEUKuM3+OeGpvij7GwS28uHczxhOeH8km/XC59L
7mGbXXnICdFBKyJdRdb3U8mjUBtKoBFdRXp2x9FUWDzrkFPJbj5h9CQdAiVTHsOx01TMA4ALmZOx
rLXdcbRgMG8m43g1g+z6dulrF1CO1dhzvA1vUisXv+3ICaqOZr7SqexDPEknf7RE1hlkvJmFGO7b
VjrTqOV2qUGal/k9SRrsUOQ7Iom+aTAMTPpxvVnuydYi8YPo58ewLIpl7DVaxjpIzXy5/NnwOUrZ
8YVOPtEKBhTU1iesANp/1/gDZSdeXjHGO5u/HAB69Ma7O6BCwk4Mw6Q6KU5hLGcIgsaUs3a2ww0i
zRjcNJ6kCfRkQE7vAx0smLwwgqJHjCXFdoe8JuCwRvz3HqO3po1QxWUny37pPvIybE0ntQVPQ0hI
JPSMTDmAB0FCRjSulIZiVYucCDedFLO834sURBsDL87vj6DiInvCel3hPba4cXdy8CqGo/QV1N7D
dod3OFi1WCtAZ4wqhQP8KyxxGP6q/qOqZc1/LW9PwCGtMqGcfm9vE/JlV/jTqotnwKpKptTSQQ0q
/8vEtit6Qy4ygp3Z+cnnPmw+2iEx09FWqExSTK2GEu+JoiASepvAaXVwkFu/Kc5//+3lJLpV+PAV
C6DM6VKIpv5cHlXga8tsGPzJal1xaabFcEQ6JkdpDECVVNUMt8Mmi1gVJZpNfv1DpAjioD+LOTzW
i3PL2Up1HUnXYqRX9/4U3bhwl09okm3MSWM7POWSY7Q4M9Z+JgMR0zP+NskK75Iy12ikgUpeqJXO
IkV6g2NVyjnscdyBrVPWsUqSgMHmvMA+9yOoMvK5sXz4/Gx9jRTNCWWnzMT5whJghysAMStHXXYW
XziAhjJajeRacEEXRlUa9sq3eSjJEUHMYgzI2etUmMC9IKORmtmMyG/exRZQeAJ1+P4TK17+aXMC
Z0LOB87Q3glTeZS3HB0z5QopKSZcZwkUATK4vaLiKJ3Ycy3wTgfTbAjyDCEGFpae2t8ZQ/Rro0yK
/mv0QSoP7uWvy+qUvYiLPjj4TBDEMPERqgIFcOZjgQw2wtxxD3oRMBxX0+EQfmBJx0dvCmIsl/0T
05vxASbOWvwvtnx2g9v/mJlb0iz/paQK42JWi25g0+P5NdBVD+8seN1KjK7QOOmv0uzSop3mZovR
GFmiXhYCVJDFRcvpDMDh02Bha/TOKzExbAUjD0pT1fh5KXHuKDCajdYp/lKJ0b7cA9r4IagFTd06
HwhbInPtSVMD2TMmPTeLX9PyXD/JDWKcnNC/x7d6oAJS+Yny9pZT+B6Sjo4+O9Vy71/GlfCT47bU
nN7MvJNx9HWNFk078zui9k4dyEzH5g+Y4hZhFuT7LKUAuhtvABQ50Oz44T3tU6B1DqI0itXRKJgf
HXt1xOR14GQM/H1LenJlCG1Xe+veLrD0Me51HkI4AJx3TX83SNC9URT09WuJqtgr1ZcjtUiutqJM
4lfRhTq+qHhKYEBwLrrDJMasl9f1f0gqiobti2pGcNnM/fuUseM09JGrN4tD5bLdfsNXxTl+kz1S
l/JWkAUWhSX+MPDW7v/D3YM56KKCy2wvnkBauupPut33Ylj8brCrFAT+b1VhSKMiq+ZPR2+CscX8
4ucHbM+U8kVZqzuhTIKo/xUlQwarTg5w7W35yyzRaxw/SC+GXLG5xE2Ub7jVPhD3D2G3oXbwOS19
eyRSOSL/OK1FQbFbZDjZJph89mDyoN1YZmuG5kYI8S6Hy6DKfe2BwvwxPa5mv8xhPvWst8f2W6Wc
hirExrrqn72ogtsTU9BV1SO3oHs3X2D+iQPgea0grUT1fDcLI/DdHz7e9EIDB3rUxRH14DVX8U5l
iamQONKddFcy4oat0/UODHrzQulL9jEoibbYw4vp5nnICYNoc6zDd2Tm+XyE0b1K1RAhkjDdb7FR
fnQLPVMFmE6Kwx43qyC2pBlmffMC1/2Ob5hw7HuFMYGUQMJ+s7ENi1CIV38DsJhAnaAv/y8HKXyY
sjGzu3qwwIiyOm29FhK7446lBIjHvI+JQUQOE9n2u2r/T3LYSi5vhoxM8QKSzjSZ7CJj8Ct1SCQq
3j1hDcJTkGwRjgEBYQ2/tKcn+yb87Y6hX2rpD3VzfOaBspruKrruDUA6oFeVeotjh3IwJSYHHniq
XBCn8poSeCvD51n5Vw4PtlTUG7YOM42KZSAS6mwxMb3rdk4Oj7U1Ys0zy06C+8kHMOaUm1VmTBnw
GIJ3vSb+Z7rI1JAhujqo7GXogrnJUaUJpyROSPlzE80pkk/tB1HePU3gIYD5u/U9tgZt06eFrcDE
iimBdolsJmisruYq6nkRy+pBohptXS5v4D3dMVpfJPn9ANKsyqlT0nM1lg+wZxPUIMnnH5zaMzNM
xWdsLNu5cAuQ1Cb/LpgYtvtbuRe7pqXxXYtlIMdOY32fcA0e7j9wsPQp/JedJQPGlYhSKmVJpY1R
XQ9YXk0bfxSde4fmnMXtydVtgFlTV/fyLfbxsjpUAQMooA/mvYMzwlBfeELnPIuqHOTE7+vaMAJM
UALkMyIYdcTPdJGkhVaSWeNDEpPNztHo6hnY9gnfylzF5dsttNxTWYOEbNODckPrl8FsjRRgO3jH
aSfapF32kvzNJMSeIN5pqQLwZ1o+p/Nw6GwoeGXWnfV3acLQI3uOuSd4EUN/wbp6fofnM4W12aiB
TAzrfGESdg43XYQjWGKy/S/EN1BQ4SvqQrZzbAA4+5CF37Wsws9zu+J1lZKDsisSdZtgOG666joC
FWUhNfrcgtPKwzQBlR33ze4A/MnOJqqnHvdHdPtB/XQMM01D525u0Xi043oYBXYmex+EqPXGRSRL
eykpWwoQzkNVfTr6oTC+IQyIdJdX6jnqo2SLrG53c5GtuYrTv+4+ztvNw7LW1n91a3k84EhsypZ4
5zkm3tWjjADqJGTEI5HI1MFupKfgWWjuESX7PC3XKACxD3uIaD72AjCzlY2VlBJ7ZBWdBOAgJ6AR
AGrSBcsI1uWpSBbLxNv4wdCZrBOonZPZMyFsbLS7RkapBSKYVs1LZIUpVVEbGGzvFXJwc4sYlBgN
lDgQybh6USvzfGLhF+pg1fACTgC4NTPL2+aVDWDCp18hEWTdI8MIvv+K4cWULIdEUkdI7ptU4Z/H
OY9lcOD+bSZdHy9XMvAP/TpIX++pSqDs6vCU/feKk/hGuKk5GYs92C9c5301iDSK7atv1aCreAeF
y6/m07ZIbk451bDgsdcSh1i2BhRbWN8lagH0gsXb070XkOpjgemz53rhQgZCPKe7D94E2zEU6gj/
mo74ER0pi6Q7Q/Y5fGYce7EB2Q5xPg5zPt8Zj01bZNpewL8JzBxkbvj3XwF+zL2MNFstZBWRtFlX
lDe3Pf7GXuUt551vev9zYw9jDwqKZi6eq5OpJx+U+3jzK2SeQEez3LiXN4/wFw5bYsifH+aVEuuX
sUg6ZbNuwHB+a4sECDfqlUozsO7WOGeQnyKBxtgQK2I/NvTJ3m7zOfDx7aD104Da+fCE3rDGKUGb
S5QGi6VPbaV9EJYtHW5Yqtm5kBiXKW9zkQU+/HizbBZIpkWCapSvD4kGCysJIj2+rM7cBOEstIGr
GqcSLN7gmKaCSduB24WBaDjKpKWv6zAOGADQdFo5VLAFk1dSAHsxgmFXJNCzbvRyfOh+rwPmr1Qa
I82ig5Dk1taDuO2z2GMLt62tC/vQjo3I6iBa4YIYGU5w8AhwqonE7oO+AEnvZjsPT5ZDl8m+aL2+
Aj0Q7DnLW1qhvZMfr1PVIf+r70jew8KaS4gfqnuztGv8ltTlfq7OHEl7XgokcDoICXmrotpvulZF
OKH4FhotHC7uXBdJCiBEiv2tJ1Gll7zec4iJOBSCN8N1Z0vZK1CnG6tqJamS+he8JcI2WgVlNy3j
7IJ7AygMVHundXdxwjDKUPA1vz7krAUmc+19U9mqpKHccM+UedHyWLXXVOGSS0q6bUZZa6jgpe0u
DMyjarOFmE9kcbQpUJUb8mhbnHpVmCoNeEw+RciEiSd27ZXbrUOycGsWnUnBSyicJXxxtbgxZixH
grqAo+nEUYXjtTJeY5+tkm896oQSjTJD3BVV68tzJRnsE3oxozM51t52glU4yvElU7VK7XXVpHZO
kGMk+4n9eZzvX5amcUBSeBKfIdSZ0Wrz9SjzPgDcpQK5UO5EEPzIMMmgi9FFecPzbffdIdt0B4oA
3DSGGB2NdqngMDgPkoMn4to+BGVIFT0xCkCwoFVKgx3ezc0wKJYg91issD6eRDCO7CbYZvlIUJH2
WE8QCtWUJeXLibre0puWhVI2G8Y4yFTJsK3UDE184RYDtsoFuAERtoPCqP+sDXCyEjpDdri1S2Et
R+x99acEtxdgbA0V31ysKnIXrI4q3/X2CTFBckSgPlGmhI5HHrgHInTFS+YtG5TUGBRo9Lb2elAs
CSz2Gjo7r07XRDWsi+Cx/PHdoinGfvt2YHUwIhVcFmGi8B1qeIC9je031eNw+/PLLbfZBiteoKJt
VKx+0ME7z2FA36fdReUZa7LR/ZJOrWs9M7/ummHJL9b8wbvCusSEsnuOYUWYpvr6J2IIR6kfg4AT
VO3YEmReI6xvGgp3MD6vTilN0kk1k3xD4pIKB+/Ht7NlREZPq55GGK5SUGdVBVl2P6VMz+crdUXa
OqDmuNYMIOYJht0NKeJlEqglHRg2qJNXQIQvIatNs3pgELYVPswwxqnOGRa3L8b2XDmyFzxK/zp3
arjlYobV5WLzDT0dzuV15ez1J0YS5ss463kxzPolCgn9Pb3olz1M9UoYAzrJl2VC+odZwOBu7laJ
ONk+DSiFmnU1QHY3YRv081l9g/KV3YVU5CllNFfAK82YQ9OnzHoybC+TXV0G29MUN75fuF06Q3Nw
FaxF/SSDnRFy8dN8Pd4Fg3VHengLmZH+UcD+Yncl5axxVbcmmYfJ6YOK8F6TYXihc1MZAVNkxGrX
ooToUE8Tost1+B5V0aRwb11qbpxdtg78ZQrLxgU9769jZXNnrGdHZWub16AylQyl5pR5Elw60PsC
vIGtD+3nSygoFrffx6sbjyrxlfhWOZimluri8HwfV4MHK5vUMXJZR8v9k4CV8JtbxIun45Hi7QAs
ZlL/MvPiUEqTMhk44fzbcAp1VGmCeoUwvQ2T9u7T9i8N7qlz6cImaOsP2MaUGkZfLizUJ+63wtQK
KvngSkg68SmOOKHn3FLzr6M+5wlbCSrnLvyQf/H/V0kh6M8Ey2F60k3mEv16RDBLenu0FJxONPGt
KJjVKxGKh5u5+JhyXsBMaGfhFB84KfqA8H8gpJieQcdd+GcbUhaEL7SwW5VkakibRw/vZ5NdlfIp
U03jqKI+Ee7EaHGYOymg2oCrA/4Ej9Q1QgsdTY27Ahp0EPr19IieNkuIppGHqTcJYhyceZiie4zz
bU96RM7EeMgS3Hg6/uuF5GWhrvSJpUWcB2hsfhCF0BWbbnghB9LFYzPP2mB4fn6I3geC0CkN5hAL
T5er5eFM36stvqSszf4+0AVl6+aN1F1V8T4WT/oaPuQ0W1py4hyv6YbnCt/+lxzEWHT3fhPBY6TX
GI84IKa8kDSX3xNhI5jLPL+YmXGU4ajPDR3++edjj19thinpn2ZJaLFuvFCQOBezK3N+T41Ko/J0
UXN9Bc+lpJmCa5N19KnCLp944Q9VogytJZ4XZJP26LZY2zR/OedI3X6CDmtCQjcRdRyO8QlWhb7H
7hFRNAFe/RWx1zEu+PqslQQLONgorf6okNvhWTIvIKj8JBLtAJvMhzCX7Fuw/MQbvUS9qiFvgl/G
EJThsSqf4msGAXTRuVI88eVg4w3R0T2RodoWOmmf6bUat0/dIaeNjeY2S2ZmFICl0vDmFWbpsfUc
PlNysiZ/zdJF9XMTujoVMj+pFeQeNTVYnUA4VzVsncmjZgw+0zjoSCD73L/zk9lNqUmY0gKzKDBV
nItn25hDgmiTx4TmawZDe89tcK4OGzJ6oLoZsNzHsUJuGi5i8KtGyINg4bWYuz2LhM3D9WSyBZTf
A6zGLxGS+/t3YIeg6GkXA27SizGR0JFE9HZQM4W6q5H9LyIzJUdIJgWIXugDISMsbQs/VEAHUNtp
GXnL8L6ZXfCMMsypWs/mLiyru++0DvuZeWaDoCuPD9ZeHkqpeemqufkCxWjXWglQvHTSI/OcQILk
p8XKPIRSTSWMKFBW+WWQ1b7Au6Qzdkv7QhlYa5EjzPW6MZxnc9b/qIcw6EPdYZ31brwkLICdZ/5C
ciY++xevmY5kVZBGyTc1Tio5W2r7dAnFQttoi+1yRAjynFQB8wBpFIE0l6liaPLjYVjmGynJoNkV
Hh0Wvn9oTR3wddwQcLdBBqcOzSvmSHxYinDM6h4DBFpLfLLkUaBK0xK5mFEi9FP6UdSMHnJTiS8K
13/P7rNR383lty0AshasLZJks17eKDhQMc+zofmkwhPLZ9mM8Nl/A1jA+cHWtzMgoZfrHlkJU/Wm
tI02EU41Dn74TIVoBy7WmZ1m6bI/6/N06OjMZclX6+m0jv8UXRRIrYspKAf8gn9Dw2ZwdwHXkJTJ
4EDScvh0oPX5BrSJuakHcTFdDKuQRU/xGovSieH0/4MhiGPMeP42DeBqd/UsnNFhwUqoaGFEUa/D
q0ofBHH0XJ6j191KcRwxYhzZL44TF98FhriEAZnLCiJeXBIC6+upQw1vX2o/ijhWyyhM87whGVih
+hRzBaHVJ8EnHKmGkMG9j2DSnrVrrxTKirDHEJLTUOggi1NYWRfJsfnTh6LusWVaqIjHx6fPVuGs
8pory7eNKXujMW6f43XwZQAOlru+U/vVan+qT6yKjOwjvCrc97elEFVR1HxZcm0qWC4mCebR87AF
gbh9p4pudiAkSV65Hqxp03VBQNrZu5goafzLqCaHLKK+rwSgiVl5RRLTgltyRd5o5Opxwd3yk7pv
BUv4dW0Z5R/BgTNuG1OMof7jyM0pjKmPObl8kOjLMisstjWEdtuGp0x/Nep8F+Isw5o71G+efFNy
IgX3FFMNGTTV9dchcsu0VkE0wmEYBD7IMWDtzf4uaDQ79kCkIn/NuDXK7TvjSu6uW7a5XyG13l5z
XMm94xjp7FhbuF17QYUsWOZo5Hqke7SdufinNctVMLxurm8PAgdkDNu0jfvmySkYR4o/P4M+AL/s
eKFGlkvhB8Qvd/8KZs9PEBpz+1Cg+QfFkVZrM22L7CEAwEmN6PxH7SgsAbHTRXhGeE9ZFgYC0vCU
G648gc2RMjnc0NdQ2H2oE5/UP+pQVRWt+CT5tK5hr3vE3cAtc3B3KuRf6iSnZybsBUnODp847AF2
m7yTULdi3my8hkrwsXz+wWzOkPtO3mtl5MCtmbmK9wCRBOUODv5b/p2Q3uYsfHnwK9xi+FLOBS93
LUHnaFaYKHYSrHO9NwvELwYMGDKMBXQ0YQfsDguzyGAM7wBQBXuik5Cau19TrWbvFM98dsYxjdPy
KoL4iapviUxUjZJKivFHly31fUyc994osHwku47BR0Aj5WjMSt0llqKIHG4DrLyltHhlQ2q0xRAJ
txL7edBDuGDkyKYGc5qH5ohuFGQovvQmcXBMqeDfDTrChIZjgD92jI6Ggj+wIq1tVbA9xsPZ9GoH
+us9/JCQAWDlchWdmY4Nqp5IXy7NCXffxiEft2S2zkintdrTM3iwJwUZYMkV8Dzfi1xAG27Od0kF
Q9xedzfStJxsLbz6xNoxQvJydYuRoRkIMlUFRM3Msc/lSQqWm+SEPo0akqwbiEwKOstDSPdQchye
qninKxTX5vDBGngzIcpRVJRonNMsp5TltBPj40rUpvf7vC2LH0DuF/TX5AfN2GNJpUPbMv2z9GWT
+QrJoqx5f+d3jubL8F7Kg0GjKFz1WX+pb3gd4soZA2H3zd6gMXt514yD7IwiLAZMjqo47LXkuake
nsFRYK/17COgXVwUzSN7yfPWXDP0S4Xdx8VITOXxcpJjn82dSS64NFeIUODLtLOZtctyNGUObShV
CPnPxrYh5yIbJsS/S1SA/DWosps/7m0yqP70ZKBsi1cZdvtaFiUgfVnt0OiJ1Z3RaImh+VGj2HKT
cmbm0YetM3TId1G3lA9xwTA6oh3Ud02r9kndG9QLtN81YJx8bsJGOWU1IrtCs753ROkmfP3jOREw
gKURUeuArRoYEH0hWTXysXclU8EMnvzgMxQVbvAw5/VGaOAV7SSxfqdwFbYPee+5/NYRk9u06eZv
sgs3gpfT4Vu+ZA5vLuJK+e2gkBfrrSjPV12alGRNusO/q85VPYkdF5910kIfYMPDOz+tFRFFknRG
NpsdTdLhrj5jP/czbqnLEfnZOeAuJsK7a37aoMXqQxjmixcJEWrKPlKccsFYSS5LsJmvfPsmwfXo
4QMl/YvKDhddQT65Hp/twzJfk+nFhjPpuhsZqxm0NfCtG3h4WNb+8vE6ZHQ9zx1u89qZ7wE1HUCo
744i5Dacag5ynW6vcWbodu1qhY3u3Khq4T8d8OO7XsY5wGyzaTct7ga/X/+a37UJv3IYCSTKoLLD
0ThUe/PwI3c8B9XVX4V/n/irnJ1dPxr1kZUHtj+yfJzyw+ej7XFvfyQiORQLTpFU/RR6LzOzyuxS
lcBwAUZH1TOsxq4LBGPUaJmVHM4gNGDnBixENY4tPqo6Scag7Sgyl5s29mUQ3tBD4Q4l/C1Qu5eB
+l7gtwXxGb+L/EFZSC0QPqorLXxSgd6XqkGkmZmsZ6ifi4CTn0JhU2B3PCy+xepo/jathsehxudZ
fSANatRoGHS085R4GvZ2aEY4WvSUiBjfCeDbP9EchrUnN6pPIVh7LCZty/SCH9ielu+DBU+S8/A4
RnRQ3YqdVwjkdA8sBQTQfEdS6M8ZmZqn3rAvVUyv3hzwYxjtjhhYldb9to5YPVJJ2mioWU+hQJ9Z
SyW5r1Jo3H6gZLOHdIUPyX0wXmWbsAsbA2Md0C2DMe9YdiE4jVr8Xs8jC3CFMZl6uphy72IrypjZ
RQ83TxaXt2tXaDTCSXEM7iKkUaniWEEjYSG6JWXslGLfoDE4E9Vv++VM2/UzUMq8If36sPVo0HP6
7G1sBtfCXG63Ie9VtFHzzILvdh53KCa91CJoZMYvA9MrbZPEMY2dIpkzzN/zT1EO//jVrzovv0w8
l3lxQTWUNfECyBic0ec1As3GGg/z95e4Lk6TrkpFJLTcOPEHMdXjxDMZ6lXBkyUJRMXOPEDoG+0V
dNpQsQKPC09GN7Ds9eYoJTRtpff2s5njWHM36oxawUoHDv2gaSvO17G5bfi4dNPDqqeBstZ400V1
RbnRWssa0ZuVFUlzMf+hbNnPU4hJagok4amBfpSp6DyBjepMm0zXmXUnMQF27QpMyPKSX8wdukqZ
ZBiY/wMckG+HKuMccUSvu1DJhvA/2EVeduHtr7wedKJTxgpnl2tmf5C9eSdBxuBZYIsL8fHeVPn0
/DkagRS7LKoycxbGNf3OXDDW2B77Mr3brOeXVzRbezNTPpZCCL9Ox7/jKOEG2VI6072JNbdgyITR
GzfWdMWCiWhm6jKtL+1WrCQgIax4+xUPFftjayMufbL3sQoZFVKrC3inH7dGsARKkUcybMrz1rsk
JDRtJ4c2DvMKVQFpGgvoexPIQkswwSuhFDChAhgtvEu9qL0nKhzK0wX+fQUxCTHiie9IPYmqS/GS
Wj57fnSvftgBS9kC7a0YsyJQRHuBgTZXY1eQrA2f8CJCtGqRJuHg+D06RVkgxXrz+1bRqVdI4v4q
HjcxBJbKaBufNrQMAvIPJyWYCfWcdIYMtecDU2dkv9MLrSeWdXM3xiJGUaLtDaArdMV9QuzMNlpu
PwnkQikwr+v62owRk933dpUueh2Iggez1FDEMCqO3PnV5RlyJajakRnR1MqxnpY1EJUWu2rewX+g
t37Uo3xYg3/lYusHsMXsM3nFZSK9AEuVNNLnt1tgbmroHN8XeLbbGkdRbJwlOt15E6VWkEPrIwtr
0iVqzcVhrtYRhDXjqGhl/c5KeW8T7//62Ntbqm4yyZz/ofv7uSZ1snOdP1EWShetRqMC0O7Jh9nO
SNTXpwDkKYjkC+JPx5Eeftt8Xd7TioamW/9ipAlErH5B/TVvJOTzYCtMHoM+ngTWKStxVfYHKR8r
cQZ5PkLbwNqw6L1zSKSAlBpgqtKPqs+178Zuf9PtYXYkKNzkeFGS7/09R3VeBj7k9rgSgbQ/pr0O
Ldhiqa2nkifV+7iEIk9v6hXr9atIMTuxG0O0qo3YFFit8kLJupJ2y+KU7rLPnSOV76pfbA72cKVx
9njNY2pN/k8OeKnZD8BVsOv625eAWYJvBoqLWnWqPMF3tWRIRK53OS5yH3ynpDv4PraDlyGxgjFF
stYv4URamDozcG12M5YMSWMJCp9N8Gr+4ijGbbVliZFWZxOt/KqVlMixGG4cpuc4wkxOpBr2p7v3
LDL7sYz0TcHjH1hRWMgnJP5UKIFuVYSaqfb2yVRcJR0DT6H+Wp7QtOnUp27aOO1R89gavgSzTloV
1oqnEoOXDmx0IsiEbX/+wOH2gIkSuQo204ye9kMIrBnxHN7lzvcV8sm1Jc+z9uzT2teG/qLP7BzL
DnTsIRArqpwcqk39RX3SVsFnMxj5IjzGsFDtvVYOyWEWJcOYH7UKeC617uFLM+H4OBRwvP7MPTXg
ImqCZQ3bOWfeNOYIVwpUucxZSbG9OCydUSjJT5lPsAWf4iXwKooWBWMvZbCYw5sm/iN91W2OkyK6
fY5fMLK9mr+o6OP5ezfDizuP0KzI6RvIGKGj2LSrx7s0EomQo3wOIZA2Kl9dNmpa3d0XXTCmI+Er
5lfqgpkfqWvXLI94ARmlwCPrKJXvijQwedQlONSXQQk2SiXOGw1lYwvyOGqdXz1eGTDRPXi+A/0P
ckVtwKfFH62h3O5gWdd8M98suBlugr8HjE+UJ0PZG6As9qcHroVJ3NsDj3OXw0JzKMo+fADUfH5h
mL1kUdDST30tWdtRYFUjA6HV87qp537NdhJx4rq5tVyWyNXpEICOPeXmDc8ObYDQzCzCIEzoWSpJ
fkM3NxpvjKYHBc3vgNg1LT53wawEVgL1h3TPgFQUspRnfcWpqkz6NbKTAstlS0F8AxhcS0hdCE8m
b3qnSsnRaUML/bA8siA8lfCNLfEA+tjDrpR3jnaFR0dl34PbUYvv1iap690PbN7L6GFEZzU4Oycl
kYlt8GF3D1yM3Ku44DtF4yYhGSdHheWZQVUKU8tOeGQ1vAeJ1vgdoW6fILE2+XPB+gTvfjMP+RFv
bXz16Ep0uDKEuKpijcTLfRXkVM1W/i+seWq4nvouAS7t4Zp6XmnjoxuR9c5KMtAyyBq6W3WNAnpF
LIsFAVwDd+fEhv8pDtwObYE3qv7fskSfCwzFgw1T9SIIh0bUu7wPaJmvQnpf/MzRl8vB+SvgCJXv
jaX+d3DlgwoBP21HfMgDAbVKmY4YZ/9Z/cBCd9LpWAmMv6asyTQTI5iWIruXpLrfKlufZvwEu9S2
9feU8cCWeVs3og8cdXiZ2HexwEAsGRJKYsGpOwz37apXzyyPl7lKXDxN2BgSpTqE4n0LKa8Ankyc
sVD0fDDgKbfdMinH3Z+3gfC3zjGorp7vCZMaPzqxWEuojNgAVgJS76dZoBJBukunBv4x2GWlMGxM
kHtYU6BH/w7Wu9PhADTY5+3CmEhJ9xG5B/+dmfOgZnLdtulmy4eq7CpgQupXjaLVi1hvWnTgDNne
xG/UffKWVB/Oq+DvtB1aWJ4mzJlid3pu2wOQTRxL+Ke2WF2O0MXCwsS7c+9+easPtQzCwFTX9hQO
aQsOJixo2KMB2szs7dQqT7i1ALGTxyIWs8FE/eHblus3G/DoV1Uefp2MF6gJIY0oIi1yHnT+OGZ9
x/z66/weV077qrxbhkFspZk8LdyIazYv9XtTYVEexOLvMnwH3IL6+lSynDNTSlOsC2Xh5Sgw51WE
nqHKeF8P2hqeieF1xd2O8W2M+WDNlbzNV2NrgBoET4aBri9PuDNx8WTHlbO5Vkxx5IJxzCV2J4xJ
zYCgb7Qr2+sMjOYTwVkSYVRYn8/3Nb8k6gnTyAySm2i7HMi56m2cXSlz9EVtuJ9FTgF+Cc0XZfZr
xs3c0rKu/n+Vvig53b1vwNa2AqKvUxCMPH+sC1li5gGBC3Wl5jjiV3+j7Y4XWXFDXIKG7R29xTh9
4NeR2THxzyotLYDgEmwUXIcZadfLYsmRaD0muIOGGjWIQxsxuh5a2cxIYyDW9VPBK68Pa76TuoCX
Dg2mplGLSwnaH7MGpRXQjIuNG/hQZSBQXdLlRg7zeHXK2WSd0lpa4OmgYhi2rdQCqQzDK1Ir/iYt
jfyLLlHnCibB0XnoksJVOxzZoAXZr9+NDX9TIspVUpf9NlTOBFvtJ7VDrqyawYEHY57abryT9Jr2
MzEr26g09nY++7cGqVWj26iMKwH/ThWbIm+CNCGpQPEjDDZCETuxzoWzh2Rb0EiZluL3xiCZmxgJ
ZXDKmXzkvRHAkD9UVp5BjFUMc7Rio7O4/nr2lWjei1T31ElIhyl6UT9m5EFLc3W079wy7HPEsaIC
nxTD9bbzZFAPFX7z3502ljkUOTvDOJKf3jpI3yt3t7giRgcRU3ZtDyJmFefcrt5LFBkg52Auutmz
dujD++UdamlDVYxkEMB5iZYuV/h9ceBVRGYC4zJm+nWUNRlHljPa64NTDixuI8YimphR96A+NfkU
5+oVYlbCQjetxunvzkApw5ThBi1vAPA4EopYDsq8RF3LUfnzcQFFlvQGqY8j7TvBJEipE+jLsjec
W9ogybT82zVZBcD7HieFEGsCz5JOTv/GVagok03x4zlHUYGFz+sTBWDDGcPTI7ow5h2XDu8vc7vb
j4i1xfh0mZ47Z8gzHnWfVaFdjxwuaunh0JXNHquqjuuQmuZhHGBfOjyPs28uPulsRe2jD61M3ADH
tj0CN5+qugqfEhKnSXYkXMrktEOFJmYt759af7DXP/OynUVOwc6dJghgk6lzlaDvwwIUOIWtzHyA
euHH7rCV/IkKt+bJ91o7F2rHoJW4n/fOP00lSeIIBnFqzTVQrm56D4m+g4Pck+mgKrP6AlbCdIdO
zIEzeVXj2v1SYHAo9IgG2Z8gJrjc6q+w+rfiSTD+1PW72Ss5iERM7Md1AIL48bFeCD82RT3omwdk
w2U2gEmxeCmDNFVl6r1MvpPaoXfjr/SerPqDNiTHOlQ9j7iznnr7oDrvpVloZuZSlFUbAhpiivHb
MWr+Gqm4xIdLoR3sX7+XFdMhLAE81J5104ix2BTKpm0HHWacn6amALLiHwUUR95KDf2JyMmsYA77
QF8PaSFjiUlFyIrgtLGG+q/8g8hFAxhZZr53UTLUppgFE4FGvaTBl1KYdAp3fOchTgPKeLIXfglC
gTQZ5AnOe1OI8sUNUoKCyNpGHIOOrr9R60otiRlhFFBfpDapkkddGKID7ZrWZ0c0oSH26mF6jEtO
fvCL62rB7eNOgsZ+cJnOtueBOB1G5s5b8UrZ4YwJJeqotyuA2Y5r8JyzWBmidBJMY40vqvXEN9HP
e/Ox03b8alElMjK7lOv5G1E83IEFGxFgERphdzIar4Kz1+zZfcj49bq/rFqAN81q6yu/q4nc/a0d
KKDHAsLwr5IRCdfubt+2dJclLU86DC+armItuCEJTS7+8c7bY3Q7d9JT8Wd3AfD/wDaDC9Bwv9eb
LNOb6h+PExaGaCoxhCRSGg+3arFUMXHvvB3NmL+y12CiBQSeKXA1Y4gyTrMCG4cTfwNVYzFJNUQY
7LG5pDVBlrPU06FicgjRiQox1GdvP6u9KrpgzU2keC315qGm4HN2XbhjoxgkqaDEl2/BzMZPZMr0
wHVKZWz+SC3tdSku3MqcuzlqkMXpSxVUe+ewxY4tgY4U9Zqb9EY9QlMRJmT0f5yLmBLkz/tujdQA
Zxb6uPNH0G2hfSDDyeHxCnLC1OGjBueGWlYIIL5w39prjCYIbeGMGTo5Lyw33SMTGfkUzbVzcTqW
diP6DvnDKzhRxnM+ZJnsb0/ixsDpil10FBrehHQWzLFbpGT91DKnTx8PeY/zMA7HxX9+GkuAmuNX
rKIVeA5gKsMzFRoYVkDSmW5V0TrVroLr5Jzx2qtKOSRbVwkBKJxoS/HhtSbMRo73SfZ8T73itsS+
cpuUUvooahK0dVCIlP7/LiijQaDJvxs1xwp3PgxQnt5KVBdEa8MwGw/H1g7XovDc26w6Ll15OarH
BKbhMPMFYi3PJ5+sJ2pD1v8hxPyKELoofBl/wet7Kq3VEdvUz+tjNWjdArIthugtnMIDl4eCtrBK
PzETmoErs3vLaiMUACF0NBWtRKXxsi0oyDuuCM+gndsMoq/1yL/2GJ2/ilkcx3cp95GsFMWHn+Wt
iDHtwOhUHGqjogQ/4jZLhN7s9Qwlg7oVy5dayI2J8fAtZDx8CTWNt+wlO9Ssk4C0p1N7y44Pg/YG
6FAnKCGitOfkFn8DqZopFSlVTv1Vtj5j+L5nHFqmpJ2H3HNp9Wkwa5G6clRHFd16lWTN6Mep1NKz
ZKs6vZkVX59+oeZ83CWVJi37PZlSwcxvGTbhuXRcI2HTUrMi+1SEZz+owjeiSpy6Tcx6rsu8ppG2
n3f2Oc6iqut0FEOQNgEdBBbpVAE//93bcwrnULtyJKZaSM4ezvdDYnQOiglyRHoDYwmxw3Pfxtcs
DygIqZZ6A/twghXpM6+tjbb+Eyuyv4qU02+0RquLXUdm8TqFSyPRMOFzniY1SEb9juXF8OnTpaDg
N/l2xDVgK/VRVOTyqy2O7UfNZz5R5DCveMyw4zWGeHwMu/HQr36WSjIiZd4SEbZPm0DKwtEgFrSx
315cKeVR4ZG81Nvlgj9f3ph3AC6fYA9J0wExn920SV0hXp28KFxm3i1pXd+J17W/M9bFxqjnaXwN
6eCpawSqFnlrjs2eDjQCJWTozh1bU4tt4tJ92oVEvJjiFlZ2PdA+ZA/UsK9IX7L1QC4HInHNez+3
68AQfCR56QoJoUmZUjPf1XOiwAFXhp0jn2S2U03TtMc2qImSEXbloGLEtjjW4xtKp9htMU6I6vHs
AnU7doz1s6C3Jk8aS5f5DXT/lHbSibkp8Iu3inNc4hrM9OYGwpzM7uFob3Q3QR7ssJNSI60LEhdO
7zvn0OHXqCxWoNiuLYAywO5URcck/Ei13J/KUCm39Ur/ejMRLUVD4IOMtWIcaAR6Xi4atgzMNlX/
sSmdS1o7uBXd/9IiLCkz9MawEUwwqCpHdmW0u92y9ewvez1B/dYH2ok3S3pW4IWogs3zieWp10F+
Yetb9a0RUtC2/1C7Buc+bQkzBXvYeX1+TKxx+zVBA3VF7EY2q44huoYNnPHc/eVGiRHXD+BwaTtr
MPRdQF7lRZ3vVYuOHOymVVC8l3BL/Uh+xmysT1/zj5uyCRoZOxbY+NI6PO3lQB9Pp/e+hUw4pqp4
2dpfscZV6XEbuQTTQ72cwQGMQZmgAz3MOLRO327OX/cwbmk3FM2LOraWySPpkyi5yYV5cAEBedUC
V9N7KHPgiIy+T4ZtnFfI5wRaPzWJKLCkKFO8y1uQ0puFB4j+CzMjlBoZ2I3RJLuZ8gWDdWQ4Rqtc
mEbEvNjToOHWk+N4D0EKv1mo9SRyUCohS+/HP/zAtJZY37cKavcDzOam+9xkzUuOOnHjG+wliWOk
0O12zRZk3o2eh2ylWZd5rjWTQuBXYzID46jo5+kw9SVsNMcQy1al9DElevz/7LIt+QoZ02u6Yoyk
mqXgym/6zYXrnANwUzNzw8FZtGkYe9BdxTkHF4dhsctfiJTR2o8yOkZnM0XImjWoKltMoN2PZ/Fb
jfm2yHm0l43G+1DLIKMqd/97I3VzA7z3MgqTLBkd4/0YUbkijv4h8XrZTHb+xWG97yMlQruRFuDZ
6wPSqleQy8b8CWzgCQEr+lwyACPLVrKzbPB/g6VAfF5KfKle0kV5jsXostlovq+7KoPSMfhhVEj1
nngE6JXJMqHhJV/bKy7quMue7Bwxq9BwQZAm/UA3PbUqysaQNFidIshwYYPSuAyP655Twg/P2f0c
P9MEWE7M6X5lUsIKQciOqT8v7rsyBTWpjjIZoz4buqdCT6kX3ocgAQTEtMhMAXM9+zs089eWcEHm
19p7Dbsxe73PcXX2k+Tmid69IQsFvfG6pul0ib4acmx5/fsttCLsRNMIFmmwFofexGMJ1f5HRyZS
aLVvylqKr64Khm/tGFOO50nSno2zTi079iXrFtovK1hYOJsqdfM5QaE8sYviFsHh5TfyG4JzdUGJ
8aoLDs6OU6WgvdCPvyJLmP+mjtzI+qFhFQa7fRhyXxaMr+4frcoSryprKtomCLRHkRBt3B6wC6I8
KTgN294tdJiu+txHa8NXXY/35OCzXvm7m5ehATblGWvtHdMsNvU7qnzEs6143CkrKdYhAVwL2Hvp
4z0eLGHs+w6IzfqiBXUiKGlACZ2YFdvDlImhUu+OXIDjIcZmcBrGG/VwUenjxQJG3KLaKw2EFLcD
CMz0sVBPfJhga2jkaBCJ4d0jJ2od2/H4uXwn3UvKJ/jxUz+4+euekDmUgTqA4sPvWt9jvVjZ0JOb
6kRxWs9NsvbkBybhqFoqkKxG5UMl3bbq6fdJJDzYEgt017xL+AXvt/eEvMn+KHbiINDkZStBe+hY
yBKy+bZecoj+YBUZVYnnbPcaTWo2cMaKfL3ccwwaFwgdK5SnJn38c+8J2vtlu4m7shIENKJAa+xW
mM0pSb5thpEuSWI2nqjzBLDzFRW7XAOToeETKRvk8QFtulVb0KXlOa7tNpyBqkfA1UsPxlXdkezj
xRp8A/rx4jhDXVyUrnmtQO/xxPA1B/2KLSebkaL1NwoQVzLCCqf1NdsBsDky85ryD2Cz4aCEz8CT
5lBDrPDC/jvty56l5Krmv2ggstpVE+3RA32Apyr/wAxm0kSgMVCFwyOFKFwp4Voq1fg2mCBqDpSk
CJPc3yI1fn7tQ1uskegPMowlftwtE2k7t4B1hjBh1ZSJyn5K41+JMgOcVGjQtWbde18eGH6hnnI8
9AOfaR55kihWwFQvoc8yHgx2aeCg3/ih27dptOzpdaBsuQ0/CGfBy0QbjaLG4jX8GsSUIuqVaPZ+
KPVa1FLZW5y2nrDixkna6Ucr+3P5NVReOFLVtzFHsLIvg21a+fuk46m+AdOUApC5B4yuw/puuMnr
Xnz1oehyhpZq4ZEwHbvoc/iEqxBGI8De5OvihoEkbwEReiaH0O32yuVlqPGMS0v1FiOIbfBma+7r
FLQNyIsBzkP3a5LGQdEXYyCt2M6yf5ld5ax2jwYW4uw2Zga450SqaN3CHfE32SnKCmP/w8B1ncTx
T8ak9VfILYfy7DO5asSzwL053bc8yPrhVydkoUMZXH+6RoPXqUGpLmaPwPCjAiKgi2ZlQTqTSj1O
Zoa2q8TgiYdH+hEiUiGwkZ+9kSD30V/vP6D8OWecfbF5KdRXQ82EX1S5ruD1d2Q5n9qLauz/+J3l
5XNWgk/avHx1wE2DVbAgZTdITSk6jT9PMfaQ9tmnVtpD4HQdRLcerPqjz0hq31pgrFgcn9bcF2j5
T0Y7B+VYIkl3g251yCxu7gxrOy0kpgfy1wtI4pmmpIef8YeCHTUy9FrNv850E1xGHwdBKkdQAJmc
S1GNcvwfE6PPdgHaWXk5w0iPRqCTLkbhnEetRJzfXqm8vND7zZky91B08Vkz32TMRC5StR9lwev3
lmPn1BmTNyYdYnk2oDyna8y7W6d05Up9MWpb6nC6ptiy1WUODs1Ilj8N4HQXUZtbsd4uAuIsFJk6
c93iZPcadvR1y0gVlw/4cGiXbmctZpvusWG51Gu556oyQgYTSPF/ZUEwaqz+rS7wXiZeyqhNawZx
9EuGeruhVahYA7KbXRlePDzseUr1f5yNF19uIjjkmHtuXn/XXjQaYbD2frAidcWTWPH4PC7R3mxy
w5LT2GUthK5G3CUZykPPMkRbBi8edn9EodpY3BLx0jcBhglaCj/bMcgd0e+e+T0eslSWUFqcwIGW
cpxLopM4wRCKsddijAgkU2A1oAAVS9GciCaGLTsOmJIzTyNMlviD4TXD1fpO3WiZMGkY1LNlqTcg
W74nwjXZdMe5GQqJKHwFs9gRALbpEU7w0uQ15JC4z7EP2hsvVELnixuhcOYTKq5QTUN4FuWbAyge
2zSuYSwEL6Ok9sdffTpqPLDHBytgamShzNj2N9+grECa/ofAmEWAHGxLJ86f3fYKWAsljnqupzXV
cTzAuP9wOkmwdFDPcTl0S4Z5m+v5lhZdAFBF7O15bXqpMp+dDpVhJF1wG7EXpUVc/cx23KLiuXuG
pkGLC8uKmBrz1trJyEY+CcSNLzk5rZH2xFPp+RtTnjhYIWtONo3+PmFAOkgmUCTh5N1X1ZAPHSm8
sXEkJ5VOSLO9yq+H4R2rvc4A7qQ4Pw7yWVphH04KwouPOFSa3r/h6RATWxCPfCPN1rG1iKys0xfC
aPlL1BmQOtcn6B+Sfn1j8k4q5WZdG8QIznx3VrVCc2I9OV+ud2xwSsNI9VQ8UB5jsEHw2aSHXZ6P
o61qG0QEXxPwEwIPmnn6EytB4WjxBqRRQxZ+IKmb0NBXd3a+M122CbhCmuFPPUifCrPx2ypXEiww
WESmAiVf1NL1qDI1Bii6miWPAEHvKlsP692i0VX0pC4FaszwFpMBWZ/814/XSADzGnF61diGW+Fq
lXmD3MUfVRRz45k3IEvh5IGzSuaGqMfq3b+Vkzyuo2J7Ufe3Of53m6/Ayp4UbiDT1Sge15OB3fTj
Y6Dx/p8KbDcPslrYp9vdw7eagFY9xEA/qft0fgubYbwb3Cqj/OOamVgcmC+rY1HLxrBxZ/7UdiqT
+9V/xGxfKTlk3vOO8fo1LcXKBp90UuloLAEM2b6L+yzLadxZG95DvRA+msEYR1aumHz8LQwDPGpg
1xuX2gaMHfzGyUl0CD8Gti+u0qZ0d06ExLSqiXoZpwWyPN53YVkT/KyWBDGIYqasKLFE9KjyjU1s
+kTgSL8aFON5McbsJ+7+N+kQ0s4n1vNV3xCDZxxpK5o33c/pQbcH1kpVvpQrjqbjQccax5bdp5Y0
5WI287ZJh5pF4GYcFf9JFPN+lgE8KqKZKoj+P8nPcDrljUOxt/t0VFGz1PvLNGMpFvbfI887sJRo
4kqpfoYsHF8r2c+ra0Fbuifq9e4Nr4jVMOwSDIvBH5KEyfRbIzEFNoE+A0Cg7UejdRsgDBm1QlNI
0X/c/GIROKIMbKIGIRj9GZUVob3S2FSpteF1v6wzl838oz4yMmENMysCS32PsmujA+DJwzbR0l44
gIIrZGn4LcfNzDUBU4ffnIJdngqaLd/fOM3Qw3VkGifVX6iFHJeymI9pUul0VDRDnnLcfaYD7AUZ
4eIa2tA7rPRq2025cGNd0kXMo23feCTpvJTytKccOGUl6ZDtxiTrz9HaH0USIxuTRQve9NPTY51o
9lwUGnYWPyqtDY+tDYq+sEvOwcGZ2cbrl/vb678/3FFVUb6oDFY+fXQ9Xmdl0ha7K4YoibF3GOC0
twg2cgZNvWdyJkfpiZTwuN3V9P9xl03ifAR830whjlDXSyCwThL/RweFhIMZLNv0VAOGm4Y6fZ2V
dvPBp8VL6a+VKXFsBm4xcS8c6GwBUgFoFrUsZYtBsqR+BRzsBEVPBVX2hLMzzoMl5I+yReLVkro5
4vmI2qlx3o5Hl2dx5zvgQqLOayOrZKmPBjasfB4JI03NSIPePO0NLJvfSKOzDZ+UMGBePFcROCFz
HMou5jLcQ0wgnMho9RrIa6d9vtqG7KkTE42cdcW3f0Y8P+myxRjBpcQN+qhfDc7jYvRicHSI00bs
ak7wTbE5kYN+MDSkFmNQsH7+PyAwZCOZHGovWqnHnl2wXfwUY3uWMHhU2/Gfyx2uVtJ63Q48W2bV
IGITh56SiaW+d7dVpa0E060Yq9hz7ov85Cs7f1GhyOnrCCnbgkR6zuXdcJh8yATl/9MOfjmg8tj0
vCWmaks8/2nHy8Pbsny4IorQcrGzkMzrdrBxXX8VG5luE0nOKd72mGJz1GZsa4GfLhEkw7PjkFsJ
hxpZl5THyLerAwUfipd8XM5BdcCTUn6IraGk3doQPiy62+WOL4u2lGxKXyyYVNq1c/p2CsaPQTPt
O0dSZx3rnOC8jUaquFiH3uKIff7Dhk3P+uW1XnkBy+mp8zBVfa9Ei6hs8lAh1wSXhPwpz7zpZZGM
t6rDqaK6+Vs9yTJNSabjKLnyJPlf5FKB9OtmzhU6LU2XkYdoTV47ZArQVSwdrT8GCV6PJw4kkjlQ
9jhgs5JCtQ3yn0/aYssOahRhl9titZ6TK0Tz0oAeSalEi/Rs/MUJ7pZL2I9o8kMZr1pN5WGcjCCG
DfdEdxj0uwq5n1wjrM4zgwXu4ef7JmBxxzBT9DaZ/BRDFcFjYb4oXYCZRascO7wSVbH5awrLPWnv
ljfKkWZb7S4/Qj0h7UaC4D9xrI8zPBlilGTyB1GocNyUJL8cqpfelUSOx0TG9tzGDdMLbqDYuqgX
WK5wmp0tlDNIhodfTLxIvmZSQ7cDTv1NaR1+bEH47ZD1jaF7Mpm4fnNHFhBE1uUDPw0Y5h1F8xHv
BQ0FlZ4HoVwbxY+q+P9APrCSTnt90EXPTDZuhoMmbdIk9Rhb78km8wRrjnKRQO+akq3AtG8oFPEL
Qg/LXDXo63KM8Adu5evsk2qYnXMw/IIVcw6lbkELCOko4K00yGf/bBGDxi9W3UavP9/9gaRjtEM0
sBED50s3HDuZfaeoBst2asXJsl/cCrR9qmGdti4CneNEBQE80avS+3SshXB+19xbp9F67nSAyuna
bXhWsKD9h7WdmNJ4M0bLc8JqYq85+vPiYU4eC417pLeG21VCWjPU22DfQPH9iFLMswHZci1M34a3
eu0puerYazUrwFj0Ykc+uY+rfF+GpNQhLK+ec2yXEOFRnM3KVJzRdLAqK3yOThEfcZOdYU0LouPj
4aLV2Dc6WV6gf8PbJLynR7EW7NjATiPN8OcY2CiQcg8+yKp6UYMiWX36OTPF9vQfoY4VhTz9EpxQ
2vEvp4+SQ9IGhIKPSdJGIriiI0wLwWSWtJsS51mmIfTpAew6ddwLxsXxut+NlWJNCxYgvjrXXH4J
CstWzBAZguaNmn3JK2o2jGODnEdBYzqRAjCHl0vxywLPosfAHHgcSZR+LlUj62JEtYjaDHSxu9cv
6zDTOQ1TQPJTwYCaqbixgu9LSG4kemAhC2Vl5E6rYZRVhtnnHV/XqeKANCDryhZeOTQASk0ZvQSo
F/lMJTL2/DqH/YTBXyRq5aJoERVg1TlH8JgMVF9giVXG2Q4etvKFw+BN1ts5iKAB3FhohoEpsrDb
qFX77UIUjayy7tuAm0DcqWQbMkTB5ayvwqPikHuJs6p/cb/fd1wdyYwv+AWObOLEh0jp1u8aNJzd
fNNNuPLGpzgEv8j7VbgMKB6BwQNGUqZf7G8XESZaFK4B0la881yHSLqey5KaPrme5lu7i2OxpF0R
sLTda5LGCxfFdMdHq3TL0cQlRLJ5QexCBMiXzt9WlZFIIK8QgKdrX8rEKYfLyuDMSOxNI9FLzWuO
PEiaJ9NwOMyK2c8HQt0ruMwCO0hQTCkGUJNS3Mle2qnQvQYCstvzjX7IxsCS2iRrzUC3L/ogKN2Q
QFHgnoRrqvSEd9o5Uw35hUFufTfY4NQ9IfpeAImBP43EcjpnLiCNlUy/Gm+qLsCQBeHNRe/Cxw4O
89RhB7hHuYucHWiRTvsaQjBnCwnbKqnMAvGIhIPNKzAwTCIGC0k8C1qpiexmDKVIZLChVCjgiDD5
m6/0alsrBKsaZZvicY/Wt5uZ8Uq2JdaIraIQgCiKe7Kbh5LDj5a+2N7AJGCLAqkuxAKUf397BorM
XFHSBfb/8Nl+dodnR3Q/ylHHK/IqXiqlxtdQfsCSMv51+CJGt8eh8PWdY9DVbpTmYrkczVLCD4I4
ckdHrYbfLajE8ZTVlTx34+14+Vkk12lC1xV/vCAvvEYAbbrSbJXNMu20qCqAfgiQ12kxKKc2CppZ
9O1atetHC8xR/MJ7iHr6i1TprDDMRHZ+3hipLP0Naz7eqglO8cgBGJPnJujmcZsTOkM+sF6dYtxh
+Igks/u7RX6+1BJtY/qeOyh/MTUnEkia7D75eshNjuXcK2yd1uMi0Gg7kXgfkmeYtlGcuVKgCNXd
5n7XXDMyR8zzU5vInm3MuHh8hm8vT+4AwNKbCx2aizvTJimclRXwW2kKU6wAJ1B52HZ9wMgp15Gt
omzgKeQdWB4ba+bD+4pTDVy/0CPVxtuHlEzzW7qROVEdjMB0B6UT2VzDMfhIZ7UvHVSKpFDbcgZ8
abnUr7+GFkzFLEaoCDmDPdWZmV2+GvBCOqIhD90K2f7rDiqTHKsbyKVViyBcdwFt/InxzOgwmdxP
/3VcjCiXg0YzgbJRzI8il55yq1WgwD6/QvNCFhnK1EO8fRCLj4ROW7OIk20jTwreSEl++uDPAMwn
wZeyTddW+4hIYcxt0NTbBQySiEERHA2V69/N5MbH7jMFJOGuTl2BUi7L6SyIZdoe5i0r2Q+BPwYj
fKgammUmUxLZ/IyeYJUqB9f1wivRRUwAV+eVBinx5UtggOC7K8KZ4vByREotetESPp/z+yUXXz1P
6PZer/EfZvaFAJRqPvLf1QNfO2pNNHbPDqmCxaO842CQASYOV8juSluhNhRZpkKahoLkJB7hI2r0
UUKa+JVG7iMwrJ7hCP0Cp6z9qYFxeeu3q1rx+VrY58/h1Dj2I3GabD/ann1dUPpT43IHuIdFtwUU
4Kl1i3VescjSWLF+66jTQfrQjOdEt9xk8HD71mMsmJUj83jxl4Ep3iRIzRnuXBAf0tF2f/I4+3Jt
gYmho+acguBN3TElN1GYd+lhGm43wVbLk/AN/rHsWv+nyyU/weWZNMguaREpAcSupW8WuTGNuFO2
dxBjgkAFTrbFEqXd0PIqlVEaUrDHHGTFqDTWxeqLVmUN7sR4F6katsbNeqqYS8Fgxs7R3VVNw7uG
MewjmFjzUIxmIgL/iBwfMWWJO7tzFh3YSZoxZEe9DnggsQnrSKRD+2b42efOBZu8ORk5/K/kw23l
8HKs5nFhaBbSXJKAljEN1Bzfnmn0DVaulta8Jpnz1o85rr19x1GRCuRACfUY+9NQAKbMnUONvIux
V/19rw2JcTJvo8Z0yWOFg576KvIOTYlsSm76PnBviUaM8k+HNggfNSf3Wrd2SFbob8UDwe70fpeu
8tSIga5lqqAyqxEkk4FJ52FjFRbW/O2hrf5ygE3LnpR8rUYGCTSa9+1jbH1jkWezF35f64ocwlJN
9tftuznUqb0bkCZIHmRqIYxsnpX/IKwVe4NKHeGTUIIoBwWZebTMoo6bjYAIIT3QoI1d0GRqFvhD
OlY5oWk6oT81MKpUihIpgsTaas4ggdeelgCRqMzmK4qfWQ/6NOOSOQpCLaxKHzJA83dFumME4FbE
H21+bwCYKR95kby59U4PGhScIaI3kEg6Nj29bOOUQmiIsM/Ye8lBRdKCy3XFqL1jds2hPXymk8dJ
cyd7ov8hHzfeMeG7O+0OrsWWBgk+dQIsI7cwd8SKJ/QD6Z347PZKnZqfZIZOb8rDBtxa0GKVkqXN
AxcEjZ0/2VC+CNIL/TvBXolW+u6Z3z+BmP3svAsSw0rld6vYm5e3KyT+Ma4VWkqhGUhoErsB1XkF
sURcUZlndeBAInrrdhtaBCypBnSzZQ0EO7ZEmxY7sGuK7Pu6mIRgGpJHVFNaJBebS2UHVpeqim48
dEoVHDB8HY8zlEVuqs6n1Lfg3LucTqQo8WQzbOSRSqrng5l8PL5iVlDJktaryKMtbrdUIqVp8N+5
AHvG9vlCRA5mJSypMOGUwldddSSQGZTNSFvyxzLjyS2Xh/7dTmWUNvoswTEPr/ivt1yb7jyZeE2a
NN66Dw2aUJe4MZMi6hF6nt0p+DRBLzMO6v6IEh7H3FXjL3B4ai+/tN3EKquaPe9zjf29zMsr1RIH
vVWZ+4ZwNQSdn6TSlorZqBwjSAbEBOvhzTNTPvWwDGG2yTRu55kokyYpngie2VOtOHE9R1caNsK5
7G37P5zwfdaML8LutzCBEh0htmtHzZg26YkXjHdvQKwASNqV1CrHlw+31GotjCVMU1dqzxhbXnkc
4cSJkkQ3EqqoiN390gM9sLX57xTP/XZs27uvXMSIBglBwO5QdS2Wd4iBdghcKhJ28fLj1JHgAMqS
4P8ZyRGtPO1gVOTzTkWVX0/mtI5k1/Do3ytovKyi1c8bKrLgKBrzGCWa9XzBveP6oGSopv89lVCp
DIoQ9O4PiO8CiO7dy8Qp9RgIdI8QAKvVLKd/05J9voXVHugpS80rDzHQiVWeYotScVG+vIsS7RXk
90IC1W+5JpSS0vfKvfsiQFPE5snpAILwi6YdPNo5G6s+YWPUPW7iodoTwKOTqSPHJFTRqb8OuJj6
jZGPhmky8ZK+nJx4KTMNSOgOkLsg2g0MZejWHjKMAbZ8teIBGx0RjI4o0xKvYssD2Iz80fK7LCQL
9FLdlBPmmu8MhJh+LLD+RePHKPsJN/EEjnek6WDUcY2RjXssqET+bridaLNPTEn/KtbSPz0YYzEi
nLeMjNGiyYCT7KxiP2ne442zeXFyx8oKt0QIeQeWejcHWE0Fn62DhJ3R8IR35ewP5DL8kWKMn2g5
ACB2gP/1lksuMvDAW7T/3TMB0N/TaH5/M4c0MmhXm67FWodg8vUlaX1CJV9Q4HWT8cV/cJhc5wbO
Z+fH3C6t0OYZ7gC09ETQPlTolqZXosUsXN2MkmOCKScu2aTU0mkQZboBsKeCz0c/pglInP6L8ugm
f+hLHF7UqovPYG3g5GQZh75M2pZr2kjJ0F8v0Awbws026e7cxsmaaYA6WHVoBb7UCY4vK0ri6p/B
G7ZeecBw4feRh/MqSUyT79wi5ospiovnYNnpCOD36a6sFXO2OlcxqQIq5QZHNePccFfLttWi58sE
3xqN9rtCY5ff3XF6ynZLQcRDFgDoKJmJoDI7+Re78C83ME42/rNvfvu3WvvMd2EYmyo+NEzCX4iA
sCYBnk3b7u5HPozvT6I4LuqQHXSm8v11oaNPq2T5lXSLHTgZK08riQq6QfTVSbbxcA6CzjNNZd4C
w9tKj0mBY34lAItxbTVZ1vRtEGeZfzfPeL1t0u4wIUMiWPRdnX7T8x2f35c6ymhPU4oaNA4FSPFg
urFg4SChRwfHCmfiW3fJwGMMU1T9L4Wu2fpZ1UexEtRN2R8/urWy1UaH2PCGLqQ+JCFErPDCQyty
b+ikxQQwcv0TwlySb8fq1s9QSL2/qPF/rI3tOrYncYIO+6bVAtI+MZSayUKxVtcfMMb2iPpFh4QQ
FGz3Qi3Byv8RUb636Aksjipl3ZV183XqqZk85BbfG5zKq7PxBHDgr1obhW5gaapHEokw6Wwoe+kF
eO/O640eEV2bA3fdtMPf3K15FJzlMc2W+WxW26TyyKf/emnXuImvusGo2S/njY05EqoDJc0HoS+Y
gB6dSR5+g6cZevDnuWfN05NtKBZdMJE4BApstFqUmy4YwtexcVGfPt13pXlHWaz8U3DOvbn/Tt64
M9khE8mh/w0V2YD2fDEybOW3c8sVWOf/j/tIbgNOOeIhCpt0SYQgIMHZTCjTaUxxViooBUBaQiJB
qd6L1UDC96u8o3A67jkhe7TXTrowTF6Nm7Tiy45AKb7mT1DMrZJR5gc6toyct44hedFKf+KTJdKF
8+sKfwGIAt9ngKbqvQjzal/l8KD2JbU+tW1qvhrqjqUtwHeY2fbxHZW7gzI3net1yPdpfaNEq198
EKckTF5Ke1Y0TC6DmwqRzWWntppl9NSeDvTzCBmHf06zBBX2Gk1MU2tNpZjgredhGxFCua+Vn8hb
e2XtBOYkQily9ilWD1Ctlny5oY/K5HO9AyGppsHRZZi85Xnapm3+/+FexNeAdzmKjFyVDLXh6APq
jI9ywtuYmFqO/a5ByAiEFOsvZB84UUnbeQ8jbnM/xrDiRaDJTpKqAHM44inlzxdsD8mOhXsQ8tDi
8l0WG9dLoqOtG9UHVOsLhmPZ5XofYl3oWsKUuGK3xl2mBK4tDpHp3KHFV3xLoAwx34Jzm7AlGH6J
xhZWLKG6TmDj6i++bHWFqdN6secRmR+LekrGtp/eOvtepjZRKu4kDhxPv9meJ7ZnVuaOhygvBLxs
LU9V3Y5IwolJGOXV8yujvufeVv1wtCapyJptyKrb8pnqWv4OvvdVvn3zpADL5pLbOPwTjspN5KYv
EiLROkPyoBsjXG7nWZIbFOL2uCCPEpp+vEZuzvQcv/gsl0sdbQo7B2Nai+wVS5pFqB8Ou7uDbSEw
EcZWU23+J/hKEb5T2dX9vdt/11IB1YH9rsHQRkBzr3q6AZGl7ebazQfteH0n0ZviWmpKS/m2QiGd
lct+g7chq9+6h9j7A9DDt6Qv92HSLYui66ZqObabbj6HEwKfqH3U/6VABCu6lJRkstU+SFWpJOi2
m/BSZZRgTJ3dsFw8fhyV7sGJLg1kastqxOVwCS8is6SNE34DtnZbkqnyLPrFGDCsN7cH6iR3XCQP
k4NWNuUIraJrqWpSHsId3o7K/8POJfDrpdYehdDY0wxtUq0ZpG0ayST+ffI4DpdZldAgt7Z2aJJR
CuZPymio20W8fAZ38KN4bnQTGzmRdbRROEE6c7T4UxYZ48YG/M9PG7CJsSpgS+ynqUl3ujx2Xhgg
dsZ98gLCPhfQt8wX82Lm5YJRQHfnAfciqG1vw3/bk7dWupFVcksBE3U5Xo+TyEMXCmJamqDKaLmX
L/kf//fIjFGm1y2RWZdmJjzzIDDG0aFVsT8lTzTrdkxQ8GvDKoau69x77O5N3aTVCvU/25k3USLl
i6QJZu/5FMLAafhjSpuvF7Z7lLmJjFS9W5m+TLnuJeIG01AXMicg1wQRCB36iZYsY47dBGnjoBAa
LCAhd7DNQx1Oo9nPTJuy3eW3HDCPadN1BZvJT2MLVATBaUcmb0Nono3SmeSTfgfpQxU6iRDOcFGq
SVeNa0hOf7u726y5n6Ms68RDrwszrrEFyEy5RmHUnHeI0fqkQJJxsJ0yz17SJbGpi1U40UyNRiCm
xwMggPrYYEX4Ofh8Rbo3h+iLhbmpjv5BBbx5kygX7F5+rqEwsFu1z4BLMluSYKIc13VM8UM0TkSI
GP3DaExV8DHHz11ECH2Fs21QUYB2++0guWrQvQTwH98eU2yYMFx73+/jcbwm8PYtAusN51NCJ3JA
boG9EffazwpjeSQJHhweSvCYj79C+SIBR6O/93vywkmf4gP0cshJHgURzulE3IGT8RRpPCm//5o6
iRlzPts+U9Nxvmj5BEakthR5i3Ku6pc2ca+Fw9fbceFagKTFn5kPtIsBYBDyoOs3lhJrNCOCvkH9
xbnH/izRi6M0hHD8co18t7DAJi0VjnscPQ8Ud3poZtSey12j1l00VSpoE6XHd2UReBRwEMC0DhQf
9bJyUmoNPYGbc1Wq7wzmX2C3tQBly78PhnnGEbW1C9axIJCwSH4PpLcjhhQrbuhHuP6HvQ2DKH/N
mVWT5TkNzSK4pinzxvEVUOyZttAaaPI48GO0Sia6txp2RBTuwlIKojb3NzuggaNeQz+nO2ZOoXYY
CQXaCxxURPTtZdxjHGckVDOtcXt0FKtm1fLVJ+zjEs9rfVal69jDR+PwPe9zY/ZC03lJuJS2pFqz
MJWx/TlyRgTObHcdWgjZtmLqQoy8qcA3LW9UxqB7ofCQQ2F+ZJU1r97F3F8yTqGAGxox7z6U5XTs
LEdjYT7ZBb7NvTlWxUfqRHIcFxsl4G8wV6BHUBRQ6xrysHK77Naj6fjbip2SpDYb/CAHLF55Cb/h
klCSMOjSKMw0p64cvYvlNbNWURjGTcurAHLn+baVxU87loN6md3QkbrZkD+TzXGBwzR/Qx9e2vC8
7zxM2pynIvNusHhQatyLbo2wbV0SZTWvEIWmS4fc5ZfNQWUGO9veFyEscRnuImAcx0yN74dqU7WC
/stLnHIWwpcal+Lw4QhZJ1UPTFePdLanZJ4aOZqhKjAnFHUsYEs45c8iTFgkM5ebt1G0s1Fkpu9G
VqlRe+Wz8hQTpUnF8FIbVvyTZKP3lT5mRW7fcH0rIogBMT50rhtFH/mN/wx5K5NRmSRhxN2KwY+l
ZpEunNqQiLMTkqFnyyClUkMoHzfPKDlgPNk3qASTqwMI3k3WHr38QmdHd8UQLwdhnRJEh118O7Xw
qtJLX1tcGnsfSX24k/L10eNMyiwBcxWly9v8udP10vLvilab2Bk8WMMOoHOuw2t2kSfVjrV/rSjq
kFwHNKF3APBCTPbZuQDwiqZtMFq6PLQK8UqnVUV5+aeT7cJcjOYP2wr3OI7a1r0ATjMrJC8fP2XY
CQDAfgjyX6a2+S2Qb6eczH9ebQ8GW6YMASbg/GbramdoGTBphZvHTvgHdsFpcGF8tgTraWqvBJjt
ili4Fo9z9F5bROeEN7no39u03q34hptCzo2W9nXvCwQGlrkXQyN8p1Pcq2HyfUsl+w3PKXBVXMRX
/oO58dCZWq4SCL4nA880NQ2DrB2uMB0saYPn5NQA3DMYxEQQluDlulfeThPXjkK/3x5ybuw6+wRN
7nwo6kNBXuZA8KZ7x2z7ElxQV+jQpl/zi4WUB/Hrtez5yCxXWGlZD7oWPGDdKLNX7Ij3MEfZUlD1
uk8BM1o8bivgtOvYku40oovJcheg2f5yaCB0dWKVa806V5QGJWi87kMai+7KG/32ZmUG/plNava2
Dsl/duaomIVoBZdQlNJgVRuOXrwW8kDusE4eFAzpJpCF6D1oekK6XctgaSoKYBVNBKPtzs2dfUUz
bdCKYkVOnXHZ4nAM8RY2oSTAKdnqtCLpM7z2plr3HWjFYoCFRXS2+4m9Rv8uVvtjfURJVlLbmaU/
Hdt8e8BuOtA2wk/eSj8fPsLjHJ3U9aEYrWX4AEUb8TULjbY=
`protect end_protected
