-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nVXCcbFVpLhJElveiz5DV0W7vr6v5f4Nk/Sawsz/NhWbl4A20LN6MwwWLsNYde2oBkR6sOopWOA3
JpDkRXC/tOzj07qi9qlkd7tk0R1kJaxgVAbp5Hp+XA3Vs1kG6RgyHcIfBoigJBKRRlpxYI3gXLMb
gbfail1maHHZQw/trQPwKjFwbvQXNh2leZ9rRBEdak88vvKzLIOMVazrM1rNfbn5QRJAEkDV/GHJ
+Mr6rOwGD+tZgJiedE8EArPWZ48vDYLH8ckIluvLAkMe+H1Bjt4EgfczrRXBzPYVqIG6sw3wFXK+
tOqQGEbUlRPnvQlNC2rUug3OJqfCguh7TT0RVA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4656)
`protect data_block
ETisSMpyOLVRoUeJQ0AU0ClOUr6jht63yAgitPWkNXigkoFYENHO3CJp24kcuiMY9uuVWVrUtpqS
60mZSMoiO/lr1GdjYer/VYQQy7KhosN1+p5jJNpUyM3fo5BmheqqNpaDsy8Ab4jo4TYBK4bBBFiV
3gJtjea/KvBU/5LM1YhS0FuoTYCSB6IFL8ZrM1B/hewHHI3mrY+7V4+njE4oY0vvpUp/Ywkold2t
vaCgAKrNshpMHTnchnRiOxCs5wy6JDsVH9gnMK+s5HgyiP48h0ETw4j/rORv1QEi4h67ZgYX4PgH
5rbFbaw0vNfLiylIVpdVPZCe5nqz5j685Hgv+S1xp1YNCdv/xNQ235uqOic9CML/vqiLaMzHicp6
7MiWAjjntDlhKYLTFYZIafazBKV9uI3qBdClrqB6UjEu4t9YrHGpNwby5tB33fQGzlzUVnyb8EV9
J5qmjTyLP2MZgirbBVtrQrjIdKF8E21H9/VXBMIN3/Qi1bko29Hm600CS8pXM5UQl+OxRt4fOXpf
4Bhhu7hsuhAHCZA/OkeKRj0Xb59iTi4J2Qhi6l4+KBB3sLES+0DwOGMHuxhA68BmTn2qH4kkQ4fR
uChesvOHCJp6D+n90hLasmq7DGlcO/zep39bk7mQ3tQBAHPeLm764q7Zrjkcr51Cm7wFKtZyv5Jh
os0B/C23eE+5xoizK60IIbe28PgzX6nZOCfw9/hdZ3H+K/l8kazqof2gq2oyxm0L6bwe62GZ0h3B
0ushJtaILNTnHjYZqVMq7RtIhaIOPl4zOM1qkWyjDWRXXp4ETN/9zoKG3Au7NSCp5wXxiKM3vkV9
PCMfv+TNzW8hIkuZbXPvrnvVnYo2az0ygM7wR0+jUc1YHiVgr9KJpzenY0eMh7ONMOwo3qOK0ste
y2vRhiGVuPd7xyn7XX7PMKbG8DiZblBbr2Ak0HhRJ0ah5RQLSi3cIanP3LoB6l2N57B06WkQ6hmc
pT4b2nTCSLRMtlz6SXm5HE4pydg9Y7fY6cqt5kY27S2NQkyRJqCboXeyAZlnpbpIdlGctbCFwi/N
kv/coovUVT8sghSXDuZY4JuPEGRZKBSOqwq6FiDPuRTCzlu6/H6EW4llu0+iTdn+TYyyrlpZ0cwh
zUOo1gtPxH/YKZFjOLuGUcnvFrHFcqz29CJDqarg6OC5FYtNweCiJkl/hwy4PsqEK9+22vzjWZjj
aazE1+gZGSb+VPudLb/m4B/LVMH3b6bxwfqhrsQghyJFr9b47tGkzXTHE3U2u9bMBY4oeIgzg6Px
OAl18e7NwHVM3vvWoCokYcsfOlQTyqVbrI5wq4WHC/q+c+QKPvFeQM5qsLNxilI9CpeEqI6x7mk2
DtqECiLUQbQUhTw9iQequ5WJgEq2bLdAHwz5cQhg6qvgV6ORIPTpFxpaTPmr03Gk+us6s1mTm2Vd
/Be8U5Mjtx5qAeTOGpcO4Iz2IeD79dPpb+nwpRnrsf1QX9erCR+nqSxtdzpnyPgmlASHjXKgPVwG
U965UkKnVG0wpZ16Cl4u4xVEZPmbm92AYQXLPoMTYYhzfHjF/d9fjwYHE+E4Q2aYuxPXHPzTUMCd
uXTEz5qLEHUlkPjm2qyPS2FjaDvOvwKHmHoJZisRY/sEcQixvDXQH6Sd+uPWk8rXqmSInq0R+VDq
X256amEagltdTZqIArPhZ4sXRg0E6Ebv8U6wlGEu1919AoaG7y/1pqpUoMgvzFfrhtAX0oL/WmuP
DK456CfhFTrARSEkuibPyqNN9aDUHddZThL8eEjc6CJ2LK1cLXjlwxZ9Ec56CIxUiFF0b0aQrJrd
QEXDZ6/Z3ts+IRldtD8T3rUM8OyYIBUIKTHeDWXLfTaxm3Zsz6vkGYGshy6iWjmHcnqsBnqKyOjC
5j/A2lVTubxTod4OJrmAEDzq2Kexou2FKFDkm4Kkpo32En3r3JqVA8Xiu6logotcuDKxiGgKzHo/
lTqeLaGW1Kx5jW4D9UjC8fU9xAEvCouXOcBup4/rqv+cNGiB9EMPmDtFZs4O1uW4M2QwJLEczl7c
i5HMKph601ScyMaI1FT7KyU6l0AJEZMHbx3+OSroKh2OeEK76a1jjANmnOyLNBWKKCKdnW9pkYNi
EhEI8FqzFIB36UuSmLXeoUH5vV4ALSmXEGQ8P5t3pkG2KWg/fqaK29mSm++ZIMvKmvpxT4OhRlxv
tHXMbpbXHchnqIfM568xIekmEzhFh3SHR0UeCdYTuQHfEOFw8p/heOFNqMagiDXaIton3KFWCY6/
9INV2kGiKhj8zVTgKewnvvWlPP594W7Lwvve/Lmbg1fob0i6+Q8LADYoyqYP0YowA6vo8m8bQArc
ELr58GHEBuvZO3swJx8p3EDrs6NYC91lAA5kfg2kAHnKYNWDShlKLyK391dyANGD5thCe4OEWplT
kqwTmCKV7ffzfRw4eO6HuVkmoersEOI1eaAkCFlXvQ56C2GuoNnvnS/+T4TynysttFyP6jy7uQVc
2ZWE06DPrKTofpNoN787fc2n0Yta7WTrLTfms3D5c0a1lZ49V2Hmc2S9Rp6WExKnD4yI4p7gZoiP
9a3v9PVgJrDUlTbcPt7DcLrzsnpQb8f+aneos4whh/AL2G2zHkWYNOSXQHAZzzwN5h7VUIf6pdf1
LJ1p23BvPb1+HgUFI0izQyKAlf3I0Tf3m1oGwByb8NxpTveFiMl5WsaNU+MDM+D88R48YKWqVJff
8BYMJwoxkSgu7nYbTJkOHLaUToNEYu6TamEI7QV9/NixYjTYYocz++IY5rod2ClqVxMsWbcCDDoy
LoalRDxJ38TXfiGRsXFsHfIgxRMFafhMtURk0+B4Ze2Vc3ms9FjtkIPczGEY2ryECyHpOPeevpzx
K6mG8y0KNEt3GzNV5soJRCr3gJ7U9tvtLw2O1xssdrmIpo/sGdEQolp82BaT5mDABdtKIWs1iFBW
hjX23dbHarIjTh1aYOXU8gcmkz7Me5CBVWF/QSpnaxViFtQ9mbB77WTks23GJ8Ak6Q+70OwaYmNv
kK35LmrnPIwle85Spnd5bXGIPu5ugLgiGzk0EOOmvCq0RoOmOoLZemZzo8C4bFi+SxiNJ5lrk1lW
GyNchSlToC5+Y+wMHT1/eemQCkQNLrQFzyPYOhjXHwC7OA5fUk28oU1WlR19iDw2GKqXhZBgRr08
R+NQWKZhAqc5Y8VAq+6e5IodbpBO22RD9yM8xc7RHsapMlOv5F+oob39zK90KCvepVnshbK7eJ//
cgY/vRuO0gucqINTplPZhKxYLh++e7xO3gTOUl0e3LP55owVoryC0uu1VLOm1+LucMAs5xCfCod5
Ynwn+PsOMbOvnJ8T1iGmouJbTJncYLD6R9BXK26uxB2859h/WsUGduGoXs6mX11l3y4qo7uaJfAf
EVrp43eUOtPrE6bjJ/+VhzuCqHVafrOpoyAXRSb8xZ4wajwRCKoErFu376v3v/LfuN7C+OEfYCtl
P6BJW7fhhg/Ojb0rMH64LIsGwCIvdyU2IaQ6X134+nfjFdx4Z2TkJ+EjBbX00NIaagfvDhG8WHFz
ZGPpiqj+FIiTNiNUtOZgS3Lq3YL8ZepHOz94EcsJUU2E95vfWRcdWoVwBYNl+ZbG/yZj3ByYGDHC
FPBfxGQay55syK+Htk7PZrayadIDFS3sK7thgkXn5tThbtjrM2YnZJfyA8ektEsyp6Yb8Q289kEC
c+QjG3w1ecXP/q/cS3RVkQNYyy4tqigBCfIC+GRZaZb78auwcgULystDADTfZdaTiqJjgpMal/H3
HI3M1wIEouBz13UZqie8QSq9TdtS6QbRCy+Xf41EoUOQ9LaAJZg9p6cU2oVXDZTtT/grsnr2k3BN
Hr6o/uNbTM+VEjJo+OscxovjIuxQ71++6+AHKyBH76amlyxDdEeLw6oBbdYX4Xx9B842dIsjf89A
1OVo7XSlQZw/adbW8A+RWIrg8ZjO/uLYTpu8969xMR1G6HWnH6tb0c95nCqiuFyEnM/PwLhjkBEo
0XpsghqhJiQXNj4iywIKlThY27sxsp4vzY4HVhsZv1fBJ7NNHr8qvTHvfohpt+lYfV6jOcy9ErEM
tEHWAQ5jgMn7IVAjTC8WjTB7mo34pGimiOKPO81UEsRcoQm9C25tLjvqBOtIi7mra7+wmEC/a/xG
ZuIGs6R8vDxUYEAtlZ9OMRcCFjJdOjdASeEm6yaRofZsS4tV0EiHBsipKXfbpVy802Q0nMFt3P5p
mGlO0t/OCzEjdiqjWBol/tJvbWD4Sm0NHlDRgXYkudpFxrUgE/9Zh5eoViqQcCe+PK6FRQ6fAZ2x
B743e8biL3kxhHbIhjStD+yp4YewcAe3ozedIqaQVcEGApsSx46VGCecY22r+/YaDm961NjQdrEC
XX+UMaR3gfaK6Ndi1Qq45W1hQr8oRqe/1Q6w/th7MYJ6zFaIHSNJtYnyVXpr5z8Sgs23E1nDkVKT
aiLSmJ0vH/jVzSDMzwmWLagfsCHNG3PFqyXGn6aqilD0/JB//1HSt5qHIWGeRZ17hNDUCyk6fRIX
rJJdvDl5kxTOgEMdx0gb8udo4V4TpnFQfgYq9AvfPWIRDrDdYpIMSMRTOZO033YGFH4A458jvyCt
861+gsq/7Uk/lac6jXVHHto1LMAxVpQl7DfTnJbyI0EshX/eD5SUk8Misz0QuPhUgczzBdQHhL/G
2cy6jASUp7uV2weSs2yNXVEFRQzu9KIeWUFNHcINeMYjUsu11U8fIpDYwkuoqorrR3fUBUgvCQz/
xDBpEN0mjazZcUbTH4YbkRI5nyC554QM8plfYXnN7TTfLVA9Ej0XkeFTY1qcdANYPgXXbX5uVLF+
Cr6cbzKmjmob+JL1bySSwi8SBGGEu5ORIrYV1JR5mQ5RQ0nOlSvcW2EvBu0s44AuaVMZ9yWO+dCn
OeOaBRU00OWlIbqrC5wVUDNvpYOnNfg30rYDRi6bnp/JHCDSyizz0Te5vuX5d5IoZogQvcWBgsZW
7OzO2MdxwOjlLRHYnPAE6opUovvada3U4P5Yq5GH4hFZ68g17QK2GhAgemKupmOZisLf2diRyus+
cfpT7QYd0y1BNG5/6qcAF3snpd6Kl6lPaiC6z6DOR69wwgEjLQm/yFe5VInMxC/yE6jJSrrrA0CD
8AmQaITmvDlc8d9qdf4gLtj396mGZ6vW32WKcv08rVuFjvHDrzLZk0WEF/fYboF6BYbhztk2/nfy
P66X7eIs5gyR7H0l+ymxLQQ1HnP3V74mmJ+EM44y+LHeUnVu6fnhXr0OgL4aAeBEAGSc/8TGXqiB
eTXaS5xynkchDb0YBpB1cLwQDSHrBzWZs+9hsuA7TXHtwq5TWL7MrqfmuCbJgHpDeJ0/D0CFwNmi
qtM0sOiZwhxpPoZvnKgrn+kcE4DqYmJSyIzCbrvxCknqJQCV+vgkYpS5mkrj4Qg1GrlPab3Zak/h
9VRBHBxsiprSTTEaJylG/Ar+6gtctgsTnSYlTpkdD3vDq2IODQjlg6KUDigP2t7ZsnL2TnSmZjnO
HghK7wgievkiBy+zl7/OGcQwN91jAnLmXjuyfHDE1vq3C3iSdfSqpj9HsfntjZw9EJktrPM0miPA
sp20/IR60komidXZrddA6+yUTVtj36BcHxQqeXJdmdW09c+AQKKsB971i5Iozxn0ZbtRZpDeO3MB
sMYqqTkNv/xcDWT0Bj8FV0IieJ4LMJiEY3fuNt2FlOFC4wHNhEVE08B7bNVj+0Sh7W5gHg9fhI1K
B80y2u2xR6oVE4JBnIM0xaNDpBJRPRlKRPLKDok/VX2Ut1Z2YvdOpR9jlDlLjMKzLDVmw74Wkb7m
M8xkEL8kx7VOZ128kT/EiDJ1E2fE+KEd+QXQ4+WlTKkoUnJF6iYOqv5Tdz1XyFcIjVqOKka7FVye
FRXe09AxltdOK/A7RdlWuH55Cy0Ih4sooG4J9WhaiR30L2vqbX/VsQjzTSKkC5DHQmlTr1MNw3nc
kDaimH/yUD0sVyzOzMLgiM0a8iS6wMp0H4eSeyU6VjseYJuS65d5OviKUPbRYn+DWMkMC7ZX340C
m8YFBpGq/CGCrgZbMpDFL82jkSnJbeBsqPzuQjGlz0teafInDo2zuDPLJON05mcp9OI4GdmQ2/N0
CsWmTCp/4t4Y+1Jfu2woCEPg9sKYU2yDQTpyUvdmAmfGu97ILTEU
`protect end_protected
