-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HtNm4bAFhDeCXynj92ZMNkP9kO0SvLyVXttoFoVsGqhgtnzQ7xcUtZyMBiy7UhDwblTbbPG+aj7F
+OVsZGzS7qiaHt+r50aOElef9fURipdzIEfL7kUuXYJMA2h85iKggVfQU5470Vz4HmyTHCUs29x2
PNmJ5fGNLm2cVpZG+9KMRMWtSnRFfSK6FOzmRleKAWrxd5+268Gn+cXkWJLgrbKetUDiqM50zcCf
RvmvlzgtYiFRhGGPuo6pF8emxtabLp85gfjbResPGwm8SbFnnHnk0sbizQq0txRK206ZTd9mXoXY
e91yC/Ki1dUpLXsg+3Lb6ctlsWsQT0ejig3qBg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5632)
`protect data_block
stKQlznaDha2U5DVf6bgXibIeBApvNXWOzgFGd5YM8f2mFSR08jeZkEbkUzttqI8JTHiRCiYuQbQ
+nf80+1UymLcuSO8t7HgjslizVrCFQmeDe8+yy/RQ4Tzfs2Ld07ajY4+shJ69EfO6f/2U08cegtr
IIoN8/an1YjVIB7NEIL3yxXO4NA740Z8h9Vg+KqMsvDyW95gTRVuzfPOQOFpc4U2dkr1BtfXxCyn
urnSicl0S8j8Ti8vG/dnVDd0ffr89gGcHgIKpGa/ZwSJHWvWXBkskSywlcJgcDQ5xtq9EoEr8hsi
zvzPtf7aRblgCbH56Z2ZT2JMuJwLY8bBEsxYDf2SaE2Otm/yImx48Pn/TwCJnWE+LXU6TbweKrZS
xiIE0XydgmLHkHBckEMgwgpdu5FoBFccMRGob+G4iRlDkoiLAp4+u5WtFLUou6Y4EFtZrgQ4atce
d1PKw5H7+noSJ3B8m/hXpNvckSX8kOAlQfqibOa6kTceTyvkGJ4ATULd67v9d0e9KKnNnsMSktKT
BcUhSzQ60bn9weVlU6KgZfMt3HQbGJQ3rUzfVlkPxp2B8WrFUgckx6qfwRYWSd76ZzweYb5SomAv
mL1CKNX1PX82P+g+6Ixc6e1ltzxsZGW+1Jo1xk/h7fzwivSSTq+hx9ZL6GDxl4JXGorRwCPSfZzt
FltCRKSUwrLsEnTgU1wJLDzzw4nSYuH9D9A1lmTaN9fiWxz/YEqBObTF9pe4B07ANPQBDB7FcdCN
K+qT+Ln1Qb13Gu5WP//xuBb4JG9A5qWJgA2llDcDVNGeZmmMCHOOPB/DAXsWgo2gX+NiTZYTbFjj
NuRZU4/VBqY+8cwlcCpKiM2p38yk+E8LDPqXyHG4QgNTN17lWkqwMZ3FlpOL26HUlli6j9DRDMDA
JyLMJUUDpRFzAC0MOlN8PkPZIUN2Y4HFlTCQtnNuwosrawORgwvVM1zmWQmiP3b25Rdn7TrsS6r0
P9+QjYjYBktE53m1L3MfdBw++aZC9+RAGJMhTKkvOQXWD1yLcEM1XtNuehHjy02qk66tT6kuZvl8
IY2qZlYaJt+UvEC+WV8Dpddq6GXTvwAyL1t3D5TCqdYcW6eGY0gosHNY9ClZlnasELZ2N1MXAq4q
vrRwJE8KdWqwNK9O82Zto72Byr6mS/9T33pkOTWEFkocGSPsgZmy3Qbr3H1yRJ2rbyruJ8YfSNYH
AuYnZIFbn07L+XUvmtBz6HDVioFr0M2XwKmQHyfJeZtJw2Bo0VVe23Q27T/Tj7iPLGioGcTMy8t+
Bg5J4HO5iaMbD4Gtz0Qyt5yRbkoCMgesL1GWjhuUelviPRAruAzcyXiSyy5841Z617Chidf8S2BP
thGQk3YunhZOSBtLVbz/hp0oYMUzosnv9NTEjjPi1dhrNlNtdbj8Wgn44wtyL7POdc3gM4BLpfik
Twd3/WwpaMhQ/uovZOqjJWSz9+354rYinTTucSqLUONvAMYSH8nLVDS40DYJvoXJOpgUDh26slhL
PlWJuH0qGFkmXYvsIlelSjHV2Fq/LvXxT/ycVMbOt+bXrGUGg9XXTr9DqaArIcHnwbIFEcvrbf4C
IVcv5LGI9xO2pWIDfLONdascRyUVO87/0rrSoRBljd/Ks7Ym1upcIVpOSeXP9gu2OCeOaFmljFP7
C8MHDObD6DOtI5N++Z81AXOae3y8aaiuC9ZrR3lb13da1u3QVQZQAaE4+H3BNVq8YWvbMImNquBG
V+uAH/6bwpPVxrEGj7WpdfXkOHHW78JKMta5fc0U3uyN2T+/lCRELxwio9PqHOybx6z8aGEAA63E
a8w8+4nq4rMTtTMrtQWFLNyjbHi7ektFPY5LypRlsHht2pQvv3IWn7F6QOW/E5w+NTegSGb5eMjO
pGKIuLFH8DAJucj5bGVjrycpOU7xw3WbjExce1HKKqxij4Xs5CyOs0hYrvsBer9YogYdHtVrhx2u
zRcBQN53BYR+g46O46jRI4Kw9IHJzedEAkeSH/o0JTJStgZMAExOb6+IG4Mu+a9d9gRGtKBAan4p
r5U51DrKsjMcQuIeOCalQzE1E6cXunPMuhFes561p+3ol+Yz4UWXN1YVuwNre+4KqxFg+4mvu3aj
MUylAVlmOKx1tiTabnUryT6i5gmlbloSo3r1G0+MCFW0rOe9wcNSfXAkFfSW/6a08IsTUu39Hy26
DfH0a+PUrTzQ6nBZVNwMuu0nSSxXEi4+Cg3/F354gRIEskvq//1rAra4nHVaUAy4BUpBbdWgeI50
kFGChDv5oyJZsenQ73N+HW258DtRRd/TY4igoNZ4RIVIdyXFre4O5C0qqBSLcc9yFL+Y25b4l9wB
BCKixuSo8bm9+urbTJ1Ugf86ME2mfKuTaaMywmHB0OgOU4STr10++w7orZhzuYD3lFsjB1ydM+am
MmwDQplD3nS9geRvQcbxi+a0ip8fVJLjL0cMwpmAzahU6oh8TkY1GMEnzef1lBZaxgGusXuqPQt3
IWlMsnmtqkEceNmkOQd8s/dC3H+I4K7lbmANEjEgSMufL+M/PSH+vKFB+UZsppwBP85h1kNvsnOJ
W8IBqpShub16NuuSuVhy9wJfTPre6lZxe0FS+pItyPRrB9oEKkYI6wA8+NPhNmfzWXg33o9pDcyY
gd8iLoJLttywFC8V1cA0Hgk8I0YWe2A0vLgBfhpyQZKvEu0ITDpgCHFOAJBWtCG8SLQkjvldaoks
FEVEoYLjwVKpXvC9ExgIDKuuWuFiwJMtokbaulVqcDtAEKiNtBin2Y9WJjXiqF6Q+S7cWxym3PwQ
DJ1vnGiUIbr48Th06KxSWiwU5+jCC5jSWGpMmwH8HeRrxTjYCZFR5xjqHguYXMO9V26B843kLb9x
0agEVe3Id73pY/OGOjLVni0IeNEtypLdr+W+DAG/gswzPPdgKmyuA+dB56ex3BJqnpWFxESpT9BC
LYWnq8VNtUOuf2xftvUNA4C5EPQ3IStm7xpbKngToxqt1v2TS3/h791bSjRiTEejS+/mFwQZuJcT
R7smzV3ms68TdYLukJLrAP2fcn5/53N0DwwJVcpHYg8xsYJt8z8RJQf7VPZhkJilavur1upmyvOz
5RyHO+jfBu4FrPT55KDgyhOUoxIrrYpRLhz52bSTWKIk9US8gmZHXAm5xjFxb16H6zmVWFiAiqCh
wJA44rIRonZEoRtcXvtslsxspf6KgqoEJkyc3XRYGS0o+mnJZCsK41MnYwZIFECz57oFq6dm/i5j
/Qby8UPDCtfDoZUJ7SDUhLgJto5370lL/R6I8GHIi+6lDNQCdiE+w9cMaDufID9DiFSgjZ6LbY+0
PBgbNNxK3BSVvqNHFFtlydxfaf3Grw9v+YFL3sybO44ECS42sHtng8F3OWY6pEdI1FjI6xJP/V55
4CvVq/PPvXab6beduY5S/CbZJXcAEQVFkgAKsgLvMXIryDpGP0px9QdyDxicomWBxEjR3rP9RRc8
evoC4mTk6VftX0E+ryvJ4nijA/S7Ct7ThDdA3fi+qfvN4HejF9uP35jEel0dXVHcKaX3lIoKFdrU
DOC2ORsF7liHKjCmr5JjYlOPQIVu+sEGVxBBENTTQ/mSmkZ/BnihfQTG1/Ef5//KXHZCz1u7emah
j1fJn08f1D2tO1rs4tSjdwofi5u9Gyp7lQEJeL4D6xPcHocPYdI7QHo68vCBHxp0K5hjDHJUrqyP
9j/dMlEZJCqjelZKbvNbyC5+GdHhMYLTVmx1AMEPpsXJd7ABCk5FG4OuwQbxBExXqrnwJ2rZ/2eg
RyY7x/SMLQMywkurTeWhMg9uhyLu4XrAOFiNpM7V0I4iZ9zBD89wq4bMv1PyT0f/91gSh6UkVEa2
6fKJSTG5jr+YBpHJHbTUfwVYVMmcCL0Gp/evqQEwHVgor8UFcrQU/H9yfQ2y8YPa2ijxtzV6mwbV
1WW7hcyzZQWSAZ9Zf0ynRBVMvEVrUgTONnpehh7qPm1hfqNYlUTdnWfjGJJLmsE2Os2I7YOj2tWW
gvBRHEt9HanAMAhKnlBZ7IUrfEdbPZmQRs2Hl5d5d5nfYTwFNYpP+chGHN3YrFJ8egHMRoSvxqS+
fxyGR3wLXJ04cey1RXIWV88kVUHdmeLdUwxlhjk9QqwDljinvYUtq7MfacElI4fyKII0Pk1h+X3J
SMB3OPd7S4jPhQWx/HHWW4VJiPUnNoYPFnJs4NQbTY042cMGUOl5BbaUf8XmFd1+rfc24SNy5RLY
QrWBGWH3lkVLNakv5e36PjApD9I5LPZYi02RFy4ryMhHMKmHpVEnnzvYe9OA3NwFh/5nK02rmcOe
KBsFi27JiFWpj/NsNo56UEov1vbJ1Jn2wvbIgwpJmAVUYq8pFgBgFVlO1KT2DANVHdYVafmy8DcE
QnaAeSXO9TprTstaJalNAiCtutYcUToq3R2ENCGEs79db4DFZfHtSEZGmPSpI8fhmnNr5hnDev1v
WrEuNTbU+h5jgoUIqlQZ0OJ17uY1rEeLeG/sT/ldfD4lNf9QiSEEGTgYMVk6csxk69YGR1BwRBLc
b514Vw1mZm9rx/b/J6eFwyOdVvrrXQJkbdIVFsFA5mXR3rLge/+1aTbqkQShmWuIt/nm4UbprAh3
z8YNAlJHNkzteviTr4ICFNq2NiqLPhGRW+UXSRniihyebe3JfW5ilsmX7HGHKdAfFZ5pH/9dm3o+
r93VtpDT8wXoV/6oM6ilC832KICSkzLV88W48GL8trq4hntA/U6LfxvWXF74gINeaK3Zlr2fKJ9R
zWaEq8zHuvq9je9oMk/Nzb7ali+d2N5NxZ40cx5IsVIFM01AbuTW6/DqKi/j0AQsV+/ZHCFCO5T3
8VT90vRqQFPRWnVPwjpc9OcO4LYOMGGgVwD26oIu86AqAq7zIeU/f52AUC5Fe5w9w4GkImvIYF3Y
8feJaF9TxA15TaYo/vKq4rKGiVye7A9uW3fqjOh8ap2jjZ+j9lE+ky56aHpULDUporYDEedK7YFh
x8PVnEbxZ22u9YzkTqkdXFZJ/TasO9ZILqDFmUDAkXyhd4HvtWxQQU9dWn9+CVkORQEyHtw7WrAa
TQk9tdDJWLvphXQ8PyMwrVutYwwvXJ6HVsr1tAjfpBvZf3HDCzHjxzLowz/mRdrZQfuxKFU2J1HL
pVFhOGnU8PwB00+HdIhIBzdouAxF7xrqVokX0JK/ZwSJNGFvsz7J87v8hwzk/1KS/BtqxobhLDN5
H5mTIRM3zdDHxvfovLT1I43thpmGcMngTUReeRVPDWh0eMsA4MTkLZOj4P6J6ILhz3LNPdJoR4mB
qfNyqyJ9aV79nG6ovtzLX0UM0jbC3pa0i8EgBUYzr1fTXNy111zCqZ/WyHGWAvsCw01e83l7hlLC
LKzvP2VJc5pUe2zVJipyFQUP7atH311ePLlAMKLyi1Tfw+vAoagJLHDg+eNsXxgP1mKTdkpZvK3V
vr+ZgBOll18UBg4dKOFzEH+8g5yl0gMasYbyDAYX0SgrJ3sID9xeveE5099DSQaZE50OMyJRWF5v
Vqpxa8uKr5vc189itcTPtxjr/I8PFrSqOwL5/Xztf3+RoTXnfINbxzB3ZzN2f2uMVT8+mJthJSWa
wdBHsl+x+FOyGofN2Af/PiUN0uL+AjuvPyUpz3OaPfRyxR8J8/ZcG+T1QY7FIlqJGtWd6Bp8ndlm
rYYp8cf+PFynKNuZQNVPt6+0h4csW8gnCn1AaVfSYv5IYT3zCNIKv3sGFrpOlREkmVV4p0an67it
yO2cQUOVHrAP2fRiNu668cnjtvxguJFr/MMF4rznF97z2iQTjgL3uD9Xq1GgbS+w4R7qrIuv6p+p
kKVE97XQJTNSKVEm+GFPvpRlrf0qLBe/T1jcgpZDPArCLAHYerIweRw0s07XH0CID7TjNsWjHnX1
Ax5eusy9afE0pNYfaY/6qlqB7z45qoZ5wCojomQb6Tz58Z150wt40g07KxFPXXggNBY87uB0b9EX
coA9zYsmYyOf4o/UjZ+aEfginqVRCPZmKE5tuNEgKYKVBiB6Gt/afOhjFivmQI0p6Iqtq25685bM
KuAuyXqxLM4IAdB1MfisAE7U9j2R3ohl/s+CKEyr4yEqwRwAhttw0i5UQtQkZ4Jhoo4gdmzw6xkc
BxHO3DmiIYjxbAvfZddYdV27VEBhSHXv5akTJ4whp9NPjRD+BM43cPp3qEDhPQGAFRC3YWwBiJiT
BVK/dUJ6Ze0rLj0X+Ni1i5T8LDrJ3XFRl2dMJ9l8LBYdUmTYNEquPYMrMZkoHD4zj0J7RvXREUim
hnLJSggcXQBTTk+AoTxdzjzLY0ZqSIgjPYN8ZBeTYWrxBQ+PfVoAdUFgt8hnOrnaHlt+Ho/14qwV
Y7a/ojYnznV4whDvaCVDARi3tXv0v868iO4RUyDXxKAIXESmluqAW2McYVqIAOjxYFON2VAaXIqc
OuWo+hsCTp3HrN7EMa8qLcqXOU+mU70W2VHwzKmIHsmzeJHkEapl1qSYAEOnoxbWT18L3/2NK+s2
xLOHJw7XsQ8wBtxCk9GDXWeSNOpYqNteQ4wyfO9UvQDsj4izRHv27HS7iKOX7VMWqpyE8vDBQpxz
Aeg8N3W49gsE7brb8Kjk1u0wOtlsu8e+z5FqQaz/PL4oXz93VA4oKwzMGxDAVb9DWX9VrVfZ6iSC
m8qUSXwiahVXbVNWVm+x7QMH9iGkJ7FHDxZ/qqKqE7uL7MiWUoYXQjE+d9Ex4lFNZd5gDuQO6PV5
1VzRJ5ghICe7Ilf8tagNp7rdqrLwK+WuC43/z42z9czf31T63Gc1L20+M/tTC3ejGsyQPvyoqw+Q
d71rGT8NcRLO+SAMpU/zy06+9BJ093xArCfli1O/CP4bxEqKjupk0J7gXy32R7kGbTOMf9E2lLuQ
GuB22p4aYA+jxyLwCW7dnQcZHVpn7h9JoD8JuBSre180JUWyGUdfkcwgpXdawgtdGEYegayG1qpm
LPcEy3p8/r37/D7jAyNNJwHk8+POaYt32HaXuoRrxIIzqrl9TIR7SIhl6QBZuhcSa90qsVlGjrv8
IXdAjlPwK8KgFC827anPoXSAWY27vXsEl/8M0C9zkK3tyuPkVO5y7Sy9LbWzeQ0cqi0NA1zoO0Wf
Educ4KZFoJdJ6qvUstw8FA21PMi+P8KVppg92gw+DxflDt7gDKJGZhePWCG0oviWo//KVlUWim+B
pe0TadvdlXT8jdnXNzBnzX6uAEOfEHAUM5/8TwcbMZ7rUocek5vZOI99eJIhdpsUHytn8U4XUuWa
55/pvIKSQ72d7JKRh0+TnSURJfCtHOW3QdbWRc7kHmhIM7eTyAboGBm0DbQsJrrNZxIurMItpnS3
uCLfOQfxlz+cUdDUbVBwA8N7pECIZI7q7qraVgYepv4LgsbaYFe+tIIMBTsJhhTPb5mlonzM1Wgy
/UMZP/sKNhMSMxfYpqI4ba67LQc14s5GYudxo/KB4jb8Vh98BL9PngDvod5F/A==
`protect end_protected
