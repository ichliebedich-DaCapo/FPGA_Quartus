-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K90h0000WYQLYDooa14xaw4wBG6NbXeZi9QK/spDdH6rjJr0UBmd0Cs1SB9cvgn0KecaS92nwz4Q
A5ofietQPivZgcJd5YWmOlLikyubTuQ36OrOPnP3G99yovptbqsJVnuLz1aQFxfQ/kadqF4WI10/
ACj8Yhz4/M6HWP36e9Gej4DNz1pEsTT7fzJIcv7qsbCdyma650hOOvpEOXGdazIt3FFucJLMIiBv
5teIMVMjXVSEh6lAb2UDXfmB9ZwFmTlgfazlHPIhb+jGWAXrQs1ExQUFGN0hQwSxqMMlL+N3r0Du
3LckQYKEm5/1mNyCESElSuzkoe+eHoCAsB5ZvA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5808)
`protect data_block
NnRc7Cc/X/QzSsLHlumuPJT/QKkZpi4AohWa5xtPGmyFgf79SOlEOp75iSW3eBe8Y1iexau47mwZ
u41oZhCD07DwOPKTkS+rWkIb9WLGwpAjdCA3MLYBTboFmKjrANmQ3loUj0DM0sPT7cjwr2Rig1MM
U1F5barduJHV1S/Jp2uQlq2ti7dHgYh9LNPkzXtSf3CMz4HwewmIXXAH+4r/zGJOUbYAVMA76L8p
BY1F2ob4i/7Atn1qvu8JrB7kYoly2Q9o26znQuS8iSwwKB2QzmEIkRVQ8ybWLsv/vRCBB7HLAucd
JVtIqVuOqrjGWmdKME7CngLCq9nLUIY79kjsmlrDI915QYa7SeyhQgC2snCvXc5dKdPUuo02qqyn
ib+OqTX1JYSLvmwGqYsULNXenNU8MPszxNHVr2lH//XtZPypNh9/kC8EsPATpf5xS48e9pI5+t86
rxfH6Fx2aqmu8FaT0RbJZRonmsLdy817oEDDsscqgxXwB2kTY2DLiGqXnxTj+0+p9MKwVUy/UXF2
PUgNgi8HscDaKxD50f3TnnI4h5I4dLz0NdF4nbdwZCr3a2d0NSwld7TNs8jlQ9KYnMa12x4qiToI
+aBbUEmmcJH3jgNSP3CAAD6RAZyAhp9fF9lSrTnyxkA/Y08shXk3dezBm5rdbzdOIM12g+FUZtbA
koslBH8n8B3VSo/kHQOiesvfqKk5O0XLF0HEfKjC66TTLesqLF7TsAOFX+psrR7r7BR1rjLvxkAJ
V4TqWiSfdRJF/AVpXD0mfmqCLhYcinJUYtbPYvJecXCp8S89n+OCrwJiOXHGEJN4ECOH53mxd+EI
z9QIohxb9Isst5MRIdbOUSbXCf/1nE4fcCwFRT7SVtKxyAinNNIHl/E64fhPnAyyw2YrISQMm4Ox
/actz0S/YzFWsm0CFEzaUpYKHzyuchkHdPY4TeyL7MuZxKKgaW9TAOP/EziN4TA7Ov4XtuoMk+8A
gGoAz+rZMuoMPtbMxnTmJWkKk6KClxFBeN+QNs2XQbUEaKHPr5Ag0dqOA+E8zBBFZtv8HQmUzfDW
jZIpPzkGozWw0RDSGXgd1IhESO8//6UZWPH6hR5uJxpHERLG1p+NDoRpV2JWOLCJjjZ73J/fgqXQ
9LeLJsdsFPBCWSNF8Cc+Lx8Vjo3255VEx6OBitWMTBpIx0zE3p5U4S8qzeUlAFlb9tRA6h3rUDGn
zcviHh+sOxZ1151DqH3T/pEvzxDYxPnZdTkKAZ3vrNTGOVpMwd9Tebyt3pFE35GK0c7HgUUYr9hM
u4dRBxYusE81iprvmFl5H5ebZ7FtyrThVG6C7zMUqXOldfG/2FubeDtkyB2Lh2yb0wHdiONxLMah
PcXvYHGLYYie4birKoBEV7CMsccHUeREupYTUP8HqVeWsvn//12RGL4TmEp4Or63hDuSKgqy3YAl
0Fs/w+HqTowCE6Qw1VGkGfwwf487nTusEtGM509Ir8dpASL8vzgDzwdaqif55otZj10Q1SAr6MxJ
pZwkcZqPFISX9KT3FoPBk1Ni8UuyP9/lA75/vDr9i3mMVJOOMsv+sYlI6WuLN9Uw/2gz/JhtjUxZ
HsYVcky7uGJlxttsFcS59Ya8tuqElNTHlZd0V+QjG46k8DKs2tlgtzH5hBOl2Pc7LV0hkCcRUUSG
+pVtXflJ0H1FNxQc3HkTvRxfFak4YYIh4bjRXfjcd0Ta1bPEUszbVWufHKw734Cql68r30iiQPzw
g0ETDfJvJBCxA3bqV8a2qTE4CFRg+AD741ajn8fqnIsSxn68cNqjihfXTHwfAXnWXVSHH8zyZfss
eVkPePayBiHO60gU6yVfW9DW86+K9wTP94abK2vTdsOD3bBzaV1a/60ImRFD5gCE/ixlVoFakT3r
I8pjj/QLAoNc+XZGDWjzCNJE+BXBvtGtNqxjdrm+OUh/txUHMfzQN8ZLOtFZlkCP6yDx0VsfGc5I
a46vP2O9nrjMg/Q3goca6QpjknMMkETlCwL2oWVX+2Y7h0NMchIKG2k0wADfZ3Rja973gWQEpCwz
fpEZINVmvuTAGrqbeF3/1hZ4fLmSP78KLth8rjjoJkxHkoMr4wBmdjmDT9HTjaYXm7tHJyed4YB0
4sKlCQKSBNY+1q0hNT/5cDiqAv3YunXN1q+bZWBahbZVHRygyavz5c/1il/SKP/xoSiwproxkymz
0iKsg4DZgT9MyOQ3A1F5yzdcXNonCUJlzqiGz0y7R3dUIfqZPGqB7lMnQ22w5ybGpUtEGeKxCaY6
WYss0prUTNCSnF0Aibnu6H97IN1rP6hWODO1J70tJwgbt5lHh8V8g3ffz5rNTQv8OKlDofxoYLWd
6BwcE9WtCs9AGOuJjhJyIcsb8cROAePL/aHXrpOPPS9I1aqzV4qBWVHK+RpWFiO2k/MxdXG+DQtp
ByF5tX9R+9QMW7sSAobrV3AXD9NI4UNOQxz03kiSz8S5+eYecy+hUtzUqDs7pWjgwzqYcmOTtrv2
iA10Wz9cA13aT7vTa85wkin/kYQmFlaNHMIlPHUCjXKUa3/eVCVZUDuB8dOrwHKCMFudDW6FBoMd
EtqpfYW3LuFv2aR+UZJnONWG8p1HBtGf4BPGriX9Z3uQD8xpjxL3p6A0UARQbNdrm8Xx3ij/vgt+
V4rsEB173xA7EKZat/orXT+64UOm0oxMvoTX4fCmDCSmy3C3iajjBA0w8VK45qu7d+MfS6gP1755
oDC7wMbiHNxnv1oaKFylcxGk+VBX4Bn8TqHGmY6HsjgVG/KYXf9esMnHYygKFMu2jDZVjX6SPEWA
QSZOJF7+DzdI6Zzz19MabEpLZ+7RMez4b634/8L2ZDliGbF2mRnviJ6r6mZmdpGZhtfPPkxb3p0I
R/f5KPAbcnfm2t1EpG76V/uXuLdVUSjGKz3IZgJ4jA8Yq6QM4rUAwGPAZ+jZBP0tRmcEJ9TZtAcN
W1foC4ESWoo9AiKjmoCrTLMk0XaaOaXyVEhc4ELLm+V5KtCJbQMPo+mhg4/CBdyFDzM+7MmoqE4O
cV7dypgBc0Ffq+fZ6mTRLMb4Kw+tfoa+bZAjDoiUmLHVboB96F5tDGqXO63Ebot93sZUAOLRp+XZ
1FcoW+AaT9oMnLKgnW3Ht2CDFoc5Zh5Fwkg/jr9Vp6G6yjxAPyF3bxffhBxucbd8yg+kJ72TepLc
rIGqjdWJe5VkFh78rKPJyXOQkhLvwuU1AfnqXaHRm7Ur2jcJrx/Ult3on5UJeboWe7q06BxxPiN6
4h93tySAWDZljE5Cnex6sL8cyY7JrQwDzUv1jsVZuIp75mFitD/1QLyYVwGM8r+0z9dM+FfWxPTA
vpwJMN5+9CWxQ56kcghAyMa3OJBvoPL0AvsLXBVMxn8ZeVIdJaYkdJRTYkoLMKHEs0qcv9UluHcC
gb6c9TV6YPivGrxszgKhISog2hE1Fo/VaQz9oek7BvMcJP8dm5RLyIPDX7k3Mcg0OOyRN0O4IsYG
ZYzRjUlCqyRV+HF7cMS3Hyg4L5SSlLF2nSC/W+ahfXeksVmOY5XpZoXP1PfBhWoQSpJGFK81korg
lcAKstI3YLRH5xA11/rCxKwRC8ISsJvLiLboVmas9oLt0eiW+nZpRrFliNDezMx2LNKozmKtmsv6
7uEtIIB9y8fwgIBWoOIXZl9zFgsTTKqP3ZdVmiF+gi8vfkFR31+UeI9O9WI7kAjN5QpehPssm0fR
1OnmY9h/yecXQ9R5svrhild/arXy0X7TycdGV4VMTqhPnDcZUyEIKCs/ha4IyHv0KZm8lDxCBLUb
hQ/5tnDkA0Hsfjfm/ySVdcX7Q1dLGFWfIpzN3MKO1Hc7oCtGdF4awN8l32+zJrbdkghZQjH0x/5p
V6ksv07mMuzd5bnnjvhmmIIzYtbrZceTfOkyA3Mnr10DtzH10tP0H53wbh9jBfFFtSkOGnyxEjRq
uX6c0EdKKPdaOJiyjGGuUrYl75nVhJ/fdBuqjt5woK1K0QhuSzNqh+PYQE3KhxoSbSMG0jvlvBoF
HqPZmi5TSpaqSRX2aa7UuQvkxBuHhblA5DTn2E1EJljISkBiU8VSymq9Ucne7m2BBF20HFRpdb2w
kmGHwT8tI3ZpxJ4ItV7coVeLignIGjKgihYNJir+kpPMQGiQ4VY9Jv9Dz2dPHl9d9EkEfvCQYK5g
D3cRmhZouF1a4dmH3jwtUC90I7GkqvRIkh1HoIHytQsxWzDD3NgeyDs5mKSqhdzPG/ZmoR8/+rc1
OMER6FuJyd1GeiSphPhO/zD2spWhmocY2ZponRWuefSO1vLpF98EhaVUcsuT0ce2WGASbHhh1HPu
gTVpe+prBVAAG2IX8HedcRWDR2rf8ibgxsIGDxMRq5IUlyHcGgH1BW+a40tv34+CTSAFzjMLjCC5
JB4fTGdZRLpf2i8fC3aldOvK5g+AC2mRWXaMJJtXYm3UAaeQ0FRq3Qtc6fcZnOhVedkW2Zsl2zfV
hN7GFWDHQdX0uxSjj0K41vh1iAc/3FTaCI9wruIHjHghLWq03e7o+O9zeQt2r+F4tiy4WDVgkEOB
65nsk/0d+4R5UUQPCAAxkyFefW/m5xS+0TtGVtGnXQIAly95q65Xe/i/hQZUxNzWiOF4xTFUAAa2
+Hf3HhE3hpiKm/ScOv8Z3/47QO42lnVr/PbdE+LjybSa5go6w5TUyeFR1WrHY/2LvbjRqsR7KkHG
26NJd+RLlTSpe1GrctDT9Yags7vvM5HPl9VOkULR6/MZH4qyX7ql2E+hzpeujgMDjgZG4Lk/V26A
bwrKREFelXaJTT1P1qfvfx9zRl53vI03ZutFKPF9qeYYvoG322hVmcVEp96pwpKYlaVdFu16Mwjp
H34yvE1F6/6ImuC7qkvAhRQIf041SfTFlyvhMcH1BDztYibwe5QuTCkngzCRPInZ8ctiCIvPgBD8
V+9f8wcrgEbJpNClt2UpsqZK4XVcjLWIBALVAJxr95EgAB2ujqPPTYsYGK9VFLRYjF8QFA5BARo/
tgIUREmGB1m9t4Ibi4B1YyqNqHeFIggA9R9bHZ1ZN1NsId3Aju9sKvUqTIZUj79BBTAN5cACzeiw
wzX4j4ka8c6HcObJFM2axNvGXhp29AAD7p/Nooq8stiLcs/F46e5oJNW+5zBdBFK+vt4Eysh4GHa
1i9wSRBvz0buvbGcT9KM/2eJFptpK71Xq632q8GQ57QKbr0lH9pZheGMhqkD+2gZExqfn6GfTqIQ
6Y5oCfaZgS/Wavu8hhj4E9kj+DuprE9GMtMCMOFvUeqdx3rNbW1boIAyfvKLS+tm7qTXHnZnLIgE
qoxVIs8/LoLh6DIfeepGmCzwH+zxv5UrueLkR4DdBXwpS+HY8Z7lEY9wCkzIHtmc1EEM2v/Db/S5
mPYwqf9hsiO+wVsxHN9NIkezPmi1LEQ1GMQlxF5tfsmkBbEIvZdcGXkgg+Jae1GXrxvx6K6i1jGl
bMA4F/FbXXEQrskFdRQpHxvC7p7PmLJA58H1mYxexjo85mC/2cJzXD+PyBeD+wlLxmK3oGIO72sM
qH561JWFCIDq32qPIq7AxBo3eP02OckPrXz9JwlBCf4jzRjVNTvYuSPIjiOhTSx3hLAl0qhR0rr9
zCJh3FyNLKh7dt0S1D+EusXKRJ5uN4tiF+nKpBSfrvBBbuyOM8BPdnsbTKzuq9qu1adNVfegHfEC
n7iIMd3H/LmqhvqjnKLMHc46ZrEE+OhyPTjLMQnpoT4x09WAEALOM8W8Dmrd+KHqgq++5wQehAkM
pqXkw9KkxkG9TMDKaRm8m1D0RLQVqMDam46R+rqbQJ5HYByRebOMMK+Yg7ZLJqTHdFo+cl4Z3NWJ
ZBJZYXEUI+He2F/tlb5P5CE9mUFSoi4GSaopData1IL66se0lTxvD+CpVY3WpObSt2GYvpvtUqAm
z6K90HV/1AdOgx4t+UHqlKO3yFWtNIo9IvmNhpJ1ekLdC+c4IHqI0xINaZQ5y3HJJNQBTBhIHgA4
HCuHKGEkiGZBrl6huq2muMYa10YTAPFoyivKLE5lxMYoE+Pbx3yPwrc/cjbZOTIOKZbKfBESIvJt
4QpgfCBNNBv1q9dq+UF+Zby92Vin9EKkMDfWDSpfbG8LS87mN4gp0cGgeGWctlHvh/FzVW09UZ0m
xAjhBgSgB4p7NJcJypUQXEsUVEcFGqZ+bpRdaV/8FZKDtW9X5soykUDlgiymVXc8IKprlszm7t/b
g/uV72xYYv+mNGGQ5ldgaHnFy/UViuYnPHq6HxcW/juW+zU2ilMGxGf2uqaQrGujWgWtRIcYf+/M
8Cmo1nZakEoFo1lRUUys89yfuQnXR1G8evOibkf4ien8hjfGU/XVI8u5ProMvBBu3P4xFe9HfO8c
3JtNQySFICCwdNGVlYZAFwwd4ftGlZFkdHeaXD+8Rw74BodlpCjIyioR7+FyAjBvrCT2+rcGl7Lu
rBb0BNXEaKCDmkTghXGL0YfcmjORj+zcw9E3h88/VQuhnuBkVkKcNkbkE4xSHsqrIn2VeaJOEVg0
Z4cR+HVIswfTqR+hBj9YXpg/ZWN34iS/m0MPgcfttswjCk/7FMiIY+KIUX7U+wYUXhHWCq6gAdQZ
/o5/7Y4/MSMZjlbVOxlXawmo7xMcIQJiY38rTfiBuFPQUOi8WKvoIh2R9M5H5TkEOjsgkeOjXibK
TyDjOj9Lzi+UKlnqd2Qyu3eRQJxfUYVH7dIusE/e5MuY+Bev21pvjFXcHovHmm/6/RwrkUHUxYmn
4cVrkluKDeCPt4o3hKmJpulEREnHKaqBsPwH7wC48gL0zJIMTVoqtOOC7JpNWfRS6izhFOhZTwSN
g0vkb59waL6OIwvRbRRy0fmeyBEogwx9+ljJiVWvSJjES+/duIe9eqPjuINTIcAXRPg5LwfCOVay
6oQsl8hPBvW5W+9SmN4+VpXMUiVSWKG5O/k2/wystYdPKyway3nCuzPVk3vDyonI941koHYoqNJS
/VwLMS4M8uDA0TLiHuaB4kt6mXgqR8wtkYe9Bgl/wTHMzEXGIPJtb5l/sEtbLzYJ1+wKTj+laoAc
yF1mhAVhMPAH1Kn4En5OaLvg30i70AS8VrgmKHlFJYbidw3u5Isyu4qyviwJaq5Qmvet0pt9sLV9
xxpokDobrVwmmuqCrdQDGsv7Nw2129omDdcTKmsK02h3tocf4n/BM/PWAaRE91IB7G9xcF4G4NHt
/9G3aGRvC9bFzDPfjEV0qVf66SY0lLDC7BmzxJBj01wPCsd8RgdsfbJ22ji1vGkgCSn7fx8pCA3U
2F/HCklHaDDcJ7AfeC+7vvG5kWxCSD2oVvGR6y0eBJO1tU/8A5mvFoLLIX0R7Vq2u/6ZFbRlBS61
p4W9WN+MutVpQGC0OudhjP3dCxEe3LleaHZIevea6r8fvTq/jlvHl7r8ZPWJ6wOtwMDp0o3grzWS
pPVyYvmAUcfYuOBn0nKZvW0CDXyNIRKqq4BG1oXXL2qq6FsISNS+eAsWmKyiG67SBR3RFbIAh8/Y
MpcJJ3XWx15yLLmwjtyGX02gJQ3OwGOc7r8sYdcUfxGORlP0B6EBj+NUNWVfzMJ8LQBUSRXwbNFT
Ne/MY6r51/+u97nGwtgrm3tQVuKHXEEtn7fnq0nxgMpX+SpuAHQgvZrbAqJaKtvcTY1XHHvui4sb
1rpbGey7c1Pw6WKOMkgHiNTxASNigcxyE03F2Y5OIw/rvsowR1lXMJgShCcc2H3Z7Cga
`protect end_protected
