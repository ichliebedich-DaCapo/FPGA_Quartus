-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hAUaH19HCRXSpGSbG/uGVsEfmE7RMLLhQ7ubhOgRK/A7JBvqXQimXdXsHxzgUTvGHpkszyUCmGku
o+bJ72LQ5TwtMpw1pm9PeJVmkAghFwFxplDlvCwP7X9WUMZ6V0ztT90aY/VVg1EGIreFSgX7NYVK
cc92ll0yhXS9vV6FCNMXJC5GTCf7Az3hpPRCQNZd/KK/51E4S8WoG00oN7mbA9L8FlextEwzK1U3
dUYuE10FxgLqaHsTHrvl6bgj1uiJw6v7qTHG049bMuaGRAR1h/Pz5RaEyU1ZGXszIani9oxVSf8v
sHmerDQH514DIeuWX/0ERkI60JdxifUlHeNexA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 44064)
`protect data_block
lPHrnQaLNO08nIN0rw3CXMhxwh3PKh7PFrw425GOt2rGaRaUv4MV2J6diz7tnjj2Soyp/WWSd3Zd
yJHX+JKlrUEHKlry3A0TQdjzi42wE36S7bh7F2EfFR5tyRWHfFCJwrPlnhWSSlRb3cX1riYlq9x+
Gwx7G8vihVDKX8qeJsFJWRNBMCOPm3LY/lQh4d1vmDUPgXYZ3rbfuzQ1sFz4Gyd3wEvoEiy9xZt2
wqztz+3sybQwpAkBYEOVwz+d7CrmsLWVZ6N7lUmUG32CV2ROspMlv/ol8611aF9OtAbso/NsNaJd
KD5P54X3VIZv46W6jFbrZkfvkGPTc4CS9INe/Id/cXd7z7TKIVFcDdGTAzK1BrP4JmBtuyqbsb+B
m0FpEv0llYKgFX1mR0Cbz/BbR5tnTZZaXZRNJHLKLEoV4G2Hr1DtFLskpvb4ASZnJ0fhydhcLAiA
MkRfvJcHJe0vKZ0DvfhBNy9eskTHieCQX0t+BH4eJOTFThH5YiKVUSEd2eCwzIzwZUDTZUAH5v4C
mVGQowmcsj3874IOc9E+DqZm8zS1NdzvQzAjGh46ykCUqNn72iuXNDSjPlIUodTGnV5Xb+pBA5Cx
314TpWMRBnYbfCg2lt9gkP3rkv8okkiNItJtdum5LDW4oQpjjElf3ZYxXa79E5rj7NN4EBaL/t+j
zWO6A+rZZ7TAKKiHCGrQ/3lnPLJhIMWeNXrIYutTB3vTjw6fjLSzqGZ4UoLkHgWaatZEYNjXGdIS
nGKrD61BlrWfAZ1j4ri6He3dn7rQi5hSP1y+2udKw8q7aTSFT4KPVqm2FgtUN14n7emIUnH9LihW
/sHfyJoXIlYa40/q+XioiI9X5T97TEJ1X/gmH0Qkmk54T4EUc7HsWnouIc5uYxH7Z9YWOyLtZnNI
pxzboO9r1S0dFh9H24a4kAIcmTjrFr+R7GW7xYABSbTPkAkqwYf1Fcr65waZwnA07Q7gwl7FHvai
NwmLSdGOglH3ERVIOnLrZdVbZH5E/urWteU5d7EtFpHgIqqyaYYNn4gCNrrchg/wzF4v6p1MC1HF
OiuVb0WP16PpmeA6IMJw+1+NMgqqqhjmB1ryk+0vyDzsTb6byYq2MG5mqtfsbxywmdx0/8oBtNqu
lql8uL5vYiG+yDvmd5fsDbED5xGxI/GPeotTc4w15+eaNDaR5JCWo6rpeuFchlspk7shHRxnBRm/
KR7IW3idEijVPwzoeQOSwsE59AraSSZsmzDE5Oh3v1u8AZOd4K0EAWc2hWfeV9y8JuaQZrRg7aqA
xfAQcsNyzaRBe0YD9M4NlC4xndjmtJJvjTVsSNlmeauED+0zTW0wAOhWDGQknsofIcB/dl4DFCkJ
TDRxf08fGUloLZGTfISSxL7YR1QPauU//6CzBz9efpWwy3qbUaDiZfr4KmqpxrL163KzbtDFjy4E
o7Jv3rbvZ9frRwvv6NUfv38XEikXBxZBE7bvFUiYaYI0Lhatt4z3enGq23X/3Ac+10QBo0kEHlfZ
HbEQMY0x+PAz1A377xnxn5KypOt5vYiKcYgbt5ZUfsxNWWqE/PP2BffIhkyRSQHEE/T3u/1x//f8
ADbP1bIA404W8itqbhVE0Grp/cxg+85MytQBQjggLEkxmapchdUrUFeScjsgVw3qloJfxMPdWOml
04gCqkg+JctV6zknBZoXs6GfWXha3o4C7zP3Y9hxv1ZjnNshgYvJnJ7itQ3l8HmA+VaXK7r8NNLa
hnr+R8CiRf/XWqKj4dCu/wwL15dwzxYfqDd/MMtln4Eyn/gYeXizPBj4e+K4OUgndry7CDw6KDGN
Xp2B7vtfrlSeAh9TLGnIkiEdmInfG7IopZo91vBswtcUjxxFuU+Ni0BCzkfm42/MAbvO4vNbABkD
gDuqqKDEqZZ217rKvizlKVxqYyjvbFiy+MRr/UvEfXknnl1jgTXQSs0cTvEdbtSrLREz5+RxN4bp
Vvqd93m4X7PCuWgVvQzJOt8OvDE+EqKjwfAqCIDFEpxH5iwFt2ewwJskG3Em93/s7VXQcR3V/XrL
P0z+L42/5c3J1AieFSiRPjA7cv5gzHrHMGshMbrJ7iAYgePpGlCpa08lShKQ/ngpmJRWepmvTKZ2
I3ULVEhuvsnauC7De3Bp6LWbSdPH6m6KZsN3qtd+qqHACCpLtqSjIWIzmlgsmnfv65Srq+pIN5rb
or5E5K+CoMITOeme8DYOOFA83BkVQiPLOqs3oWRaBaC/4I8x0Z8XpMCinCIERtY/9NLNoz+J+ys4
k1AQzQHeEtigVLp74D9pY4Zau/rOXaNK59SU2DEc8w3k6Xn9OOvx+MTxbAc38eOvyIyiMRkRUm9+
wvRE+TfbKcsw9VQnh0RU9Y4YUVcZgPBkAnsgsQIZFsdTyic/0gJ4oLPBbM6S8SMGy+rFHa5AQnR3
W6en3Nigi1bQcy7ka9tHf66QrO6mzpzgnQjL+1oS7ZyUJ7iR3pP6epE1yroqXxJFGfCySNfM8dD5
4K6l1JrJGlncQuwBEZhG5u8TYS0xtSRHPU9ux7D+LJUwkExyPaIrfpr3oP5Qw4MkFvPsugwjb5F1
+0RhUWlo7NtpPhPQnUao5xvQ2eOy8yZHbVMzBbfhA1s7s0Of/ue84BusXa1JJOeFGSjDmiFw0GJc
ROy1Ts9zc3b6NNidvsolNwqxRo4Ua+wUlD5dKDIx3x65Sj5bioxEpcDo76U6G3L9NyU/EU6qC6X3
GyFReEY8rFB5AIMxSZ3e+g4/0DOwULFVkxUl8C27hlaF4iblbb6GucwITYufWOnRTaBYRHl96+3L
m2zSU9lD08r6aZeG19He8amDm7IrbYWtQa5XH/wCJsfxF4QWbgIT8suVBeMXxz6ZLLkHDsLSbkhs
LaFOYMGeNrBj7O12a1rUP62QW/wqArSawOQxSOwWtjfFErFjT055cxOQTWopG80RROob+/f+RKRZ
lOFpCHs/KJ3WD52e3tdAhO7PiNTZxTIQXnxJMPAwFl8vldVLHQ7YfKxuFpDse8qkiJcHtIRckPJG
FAei7Cc3n7XYKZVn6xL2RAs7DqfY0tJuhAvk28xRdhvzaAnDHVmJf7bFx4JrXjdePeyn+axUDd6p
1t+95mVJYWoA8Rou77vF+jGSTju/1epsGJ8fzktLgjk+xSACG2ic82xha6hZq2IEUs77OkwwPXJq
K75z6tWdh4/u1jow7PfpjILZl2g1j2VEeqUwVVffkoxNhxWhbdpKP6M9EM76iNn4VOAji8h/42Zo
HFDzyuaTk4YhGY/aSJsFmkm8vz7HxKUsD0M/zCBGTGTNzujHPLhoR3RHjBw/leJhPa5AF17mKTRr
qzn0pvlIigONNkOiUvXH9RVtCJtnye80K+H6rPcqIabGBLcnz6cTt1HkMN/nhy/cvIv/+fdNjDfD
lZQsI8i1jVMH8TARfFVaCuHFv8zmR2ASbjgQDAn+LS55sVytnB15saDnQc/HP8vwUZyKZxfDwi1o
XXzEPivUxlx4SqUCf2KOi0eY3olmjAxluoXynOh/9I3gCBkSBFW8LG/lDG9DUfmjmTJaE4S+R1sO
ujzDZaMOww6ko2ZUMipTZqueskjGf2OKKL831l53Xn5gbPw1bApHEkW4WZWWNn/8hA5D31ZgS+0p
l9p8vUoF0hyRlvxLLoht5TcKJvSdPy3Uulh8eHgd2UxuXhyPnoHIt1wmYJxTWszkFBp0pmsZzhVc
yZIIjl+eJjfv8sB2vBlHtVsmnmx6LD9q1mytIDF+piCoFdTumOlA7KnLQSilaF4+JW8TyGlCFIry
yjjpp5NTwIQ6byGYA0+Lz3sI8WdRHL4Uje4va6GesVQIQiau1T13wbf1qcXvsBqpGeC8mlMfU2Xq
c7VerFMRdCXXs7g0clG2NwslREwFv6b9WLn01WoFG0YMSyGKFmpX/65JutnrvVcuqohMxrUhDay/
mqUt6gc7hDkYpXQ7/BSg31AV9IlQ3SG7/+jN+2f/ipZOR4SgupXxNRMUPEutb7n2BltEhAFuAXCt
hMliDW+X8AbhtR3JXWJs3yIWRWCg6K6es1qTglko8wZZpi0Cy0h1RVbDxSh6SVKqe08WwhtPJ4gR
mBXaTp0xw6Sx4cIb289EUf0jIXMM86wT/qE3V6CE5peYRqa420oJSgrcrzhMppJcR7C14woM+hvk
X45zlNp7Wb8OQq2Bk4O5qfUX7RJ8kNa8b8pjIHKkHSW4avdxH1M8agljBFvZ5fwcIEWUBS/+QUiv
L2yykl76xO8596PJs3ql9fxBEHaS0pF4Kakpm2ZX2SVNGVGNj1WdBLKGAnMp5aKE/B8NijQQWriU
bvvWrzR2TB1rAFVBdRNXBaq5OVdQ/M/nczo/irBqcwHechjANLiGlfShWe2lq1rHmdst+RVD7dC+
J24E4Ua7Y/Ecla3hkpYH/NDG3U48SC8HB1hsfuXjThlNmGe7hySnv6i+lrg8uiLel0XI51RczaXB
FUz/A6dSlKhIOVDAs4pB67uxaxbqFh4OBWZLunbPPQp1ya0qpQzEMR56evseFUCe8Hlk2wdcE4Ds
tG6nNQ6k0lY9w5e1KzKLf4hmE5yLvDHsw35/RQuqXQJK4KMpf7HVhYR12ma7L68VHjQHg6v8JDe7
XQXESO4mcEEQPt9WTahApEMYX4mlDKZri7vZjJM5f9qOcXfN1d6Gtg4OBGjjhJ5U5rzF30N4iUy+
1w+DkSi9Jcj+MrY77cvWRc3rtOQRpOQmfgei6cuL+EF43vehqNZ9SFkh98As8o9GDJVI/SBZz+oO
jfdRXui9sqI39i8Cf+zQVstdzTSctSy4DoRYFjwxO03WvNz1iTziqNK0DhsDG6/qSShYj3d1gxMc
F00VVgj8yQUePJhtBtFh0llAJkuSY1AGAxskC4WyTArzGn63vdSB3sWl/f21OUP4qGaQWgBZe12e
4cDKaHHHVDUZ68keG5FSvMGofG6Nj5ZxnHk+riV/nVYnS/qg6sKuuLigSVgihqVByhs5eeW2Evax
w0cDSHGrN8N4fvomGFUk8aPmeDkKRSy9GHTk5XcKBRhSTxJxS952Ne3DWEUfuROEc9L1dx5ktwo3
kwxCsvHceuvPp/6WXLKXHd+SXOiaTcDP2uSUyzcvzMzE16JhTLd3KdtqjHnB0FHnR+qghQNY+qXB
yAeNvtLG4Z0bTE9Gk5Mkc320Ve1RQXazz4uZx53N2RwdzzGe4uf4gwBBcvSsQePcb9A6NX6osaU4
7XYTqRlU+pe20m5XlEMCj9RN7aQSydLtclLRBW+q83fDZ3FX4ErLHSlzZbuypIa8WkS4Ldurq7Sv
rjOLRMOcMR0EqdVeZYOFjy6es2Ojpc9Hwjokpx4ynv+hVytnLMLXz0T47SnhtdSJW9IJPicAFKWt
p/SjhxEy8MlJVmq/CykJ9ohRSvETurDo/D5CMsvDNiBssR6jCgMoR9sP7jTHWZr3IpwVh3C3bgZU
vx6lgv8fV/ATr0sl1T8KGsj9a1Uw+lSfRpYsWnjXo4/SZE2RNMt6ks8INGxJTKnQTma6vzQlN336
NQcyVzuchlCbHMKK0XE1vSunq3R/CZc4nx8epAa0uz4vbnLpJoNCz9iMXoCJ84tWrUz9DW2Fx+MK
QQked2dqsQ3xmhRjuNGaDWRBfv+efrKUUyQZQzvCC74wMkz58fO4IY8iQpUSdhnN0lkdyQIuuN9E
9EGIrr936PEEjP8yclROjm/Nh1SFAv24mneCHUdZEGOxCPHHIT2VaJAhxX47jr8gfOyUMf0mvbjZ
gQ3AyS8JeK5nBbBL8zzNt2k7G9mIqJj+hgsB/Md+DE2JZ7Wd/yyu08gpFFM6NA9xSaiG7nP//zMI
AGt+uIif2jrwwM44k6kj3y4tkZwElgPRLrCHOehEdibByr+Xy/KnZHA5DxrVQjm94q9BcseXBTeP
s5uaLW95ric4c5i7hCZRgXerDxGetKzfZUw30l932+e57t4UBXMkCo7vAhophRW31rXtfKBkeGI4
7gpKjOL1ctHV9k7YMSIVPKK57rok7NfUgIPuJezvBsR3hMMRspiEszg3yqrJNU/oVkm2qlSgvmTH
/QPCXJUQo3ikw7Ewlvj9TxmJ0AOGJS5If2HmWFAOMDvQFyBsc+Wc1XeBnXSG9zw/fuXO0kVW4TNg
z/0gi+JghQvm76j6vsKMCgUwjgqez0+Akq1xKPikHJTjYGvXXBctjmyGgvojeH3zESuLL16obknE
4wGv2xpDAqPZFvIkr0Qqx92LnbYmMtUQNRS3zXKvR2+OpFxqWZhmmnORUs8D8Tsurqo60BgVo00d
pAXEeBgSlKlK1wsERCuj71WCRfe38CyfRq0oYAYfDneelkyQphwW0ok7sw87cljT1lowdDOMsQQ3
Xb7INEZZi4+nc5IDJHZ0hrYr+x3SDFeiSXSXiJ0Oe6FXRsjK80GAAgZw8YAITxv02/0csv1zPLBO
K+X3pcgMrEozdWV/GoHZmTVWdDoptsroLk0pxNKgX5Ee+WM+DtYRbZWRTbHcNLA+9a7AMfmRWZIH
zS+GK67Yw5nWW2L52T8xVw56ye179zxGsxjfm6Jbskoqj5a6ZriFeQgQKxPS7GLK3/XuMSNRvC3u
7mr/7XIQAuJ7ld3KND6BWBof8ljqNyM2IFxPidt2FI02ZP6RvjAaffEwaS0ofN1VkS/u3835i9Vo
2l2QSiMueK0mI5bUjUP8gmNTKRpgPNKYfO8WPJuuZrANYabUeZ0aeUoR+NSR7Yjw0qINuTo7eV5B
PX7RNlkZoUXsTefJSSZsely8TZDY0Z72k5jI3eAqeRBqNAYCVAzpaJtDPRAN2LhbtHpZyDFgzA2W
6LLf/7YUXZnGKVI+ggzAzm0OggxypLA1Cco1I1cPIGJznJb4zcCmqw1fE0TQQFbuskvc9EJWHEgO
ucffgJ660I9bRGLabO4CqhsfusAMuqgrnGt4nB40xDEnoqxlbhFNoLaEcwhLUSdijh+YS0dNV4Lo
ZBoO3bbAwGMgqDGHg9i+z1tMmqIh5qxULuJILn+C5Smyn/Jgi8wgD0KUtXhFCnmDNuLw0HNZQPcl
QKRF63nR0ahWOKx9CTyEncutnMatfKPT/gl66qtCysTIL7t+7oF/O0fT0dVX55uXM7bSF5xl+3pu
urtDQm1mIFoIv/nibrQ5mwJYbgZ7IOTXn1ipmySF2PcbXsT4ld9CRIIzZ+TPmMFZpU8hGUPA5mVT
i2F5yhVkXkP7qbLcV1D26lsrCnPHEfGiCUZwRZQLGOvPFPg3oiJANjW7kfNBkCcY8AkLyqaG1vTw
Zt3JrWP8U8o7Xs7PVeP44j4fYY11Jj6gdDyA+quErG0mQAiQOSF+9cTSdBinH6yPeo/2u1VXliQq
Btx326L8D4C6yJCF/hQ7fSkhmyi7KptEUthql8pJgjB1xMzYw6nEXbf+0qd/AdKNSaocTdZBuos9
IjCvxAOt2HgKworO3WtAKTlkSHHmEaWHqvhAOR4uykiwp2oQ8V3EFim/xLpmEL9MC4Qt4hlV3XEA
QwEx+qCEes1EjstmFmdHDVtHI9mTsJCLj31tIy9z0gBL2B90Gyg5hIOIz+0C2zbreboOQdMDVgMu
akanPH40avhTqDY3XBEZpUKwr+eO2bim7jwnAo/D4HWvKVzOP16bju5A15cJxaB9QFMV/yjHcmgr
w6Exrqa5UnX/qAJohYhvkYk8ZCGsYlWeWgabTYT9FO7Z7p/BnhHEC/AzkQLc1cQcXnHluILXwrlD
gHkonqcFkNde7w7wSQt8jUEQsaJhEVozElYIK4wzuqT3BVh9gGJJIU2pNl1gaUvRbmVIJ2JQ+An/
rs+WswxvyGQ8jR6my4OxVFhxFWEReKkffSG12c4FYMx8kLHAs8fUWrwjKgjrf2w4F0hxmq+9fi1E
h0hkomPUKfJvMu/ZC+YN/DVd5CnV7WkSoqI69SVomi+WNapJIb58nZuo+5Tl/Ky5ck5Y+WBv2fu6
2zrzDXOQZHJcBsq4+s51suEfBPgyBF3JBddLUGMQ+ZNIEsU9HFJH5rfFZdMSpoG23fL3TlXxM+4i
s8QJQ6O9p7RludRJOCIJQl04VjhCp1jfUllmizvNASIbBRuLrzsOBgd9A8VC3E26KONWVDf+ym7F
3Iw2ogIzxo/6G0LvJKwntAQdLxUXBJddQiUrsyy6tgLOH8j6V0VJ5TGfK4BiKqLkpJqMcAmdbxL1
QGkkkqWrCXs3A1Lby2Qt83YTREZnTNO8Yqe+UX26+IFrK0WUnoaE98m0z4hN70WCfZ+UIvPQ/pYk
D7Wiv0WvseNhpXXigOVk7wKTNXqjKXgJ39JhrMS/tGX3M6hBs/I7YanKXlHIfM1IwtCOpDmSmyCq
JF5THTWNrIqmeLIuduhsS0ruI7+JjJrQMmKwmqHgmdIzqA03dhwcL1gXa+O8LHjCmcMDot40318C
k+n25MrQhiMeeDChltQoYl2+7sWCFDtxYKM73tPRGXjJ0qmOJvwcXXP1DUH2e1oVqP0ox1ruoBBr
vooEdEh40TE+iA/YCJ0KJCbvvOnLzxMrxuluNA5LlKpdvHi1J0h3+uF3v6Urjw1fjEaH9RokWd0K
PaeLnwJLd/afX2jtQvs/GrmGR9mbGgHkY+XuYvS42+zXHKg3oo+jImagZ1ZprWBS9BI+XIPzTK0p
r2MxX9JGMKTuM8p4+nOvHwJhIO0+UBMb4XZnn9sOifZYBkiFIYtjo02UYAti/R5TaI7vPb7EZQwc
oTA0FFShNNQ7NfvBRALslbfsYx7i/yzeyuv7KSvGZqyu4VHtmJRgsS3WYBz8TvttocRT0qWaoMQ2
f7YUM9DcidnSZDakRHsIHxjkhM9vhxqpfqkhCWnFtBojZtrR556h2l9TW5duCFwlAg0oekJYfTQA
pu1HYwNrbgVd+DZSC6kOZYBdpTIOjAToQPn9LIFpXTD7ikk3VEpbXfp+E+LEiL7CpEGAy/l2OYO6
RDE9Eeubc0Hm2Eg2lJHwfPgBKzc9FsfAUhOUF9bAETt6dHfitcJ6IbXJEpWjT5YpMihE3H7Gh/Gd
lTEWWDO+yIvJgdNUPYiYnBR7/dA1hFE0lNlEOC+fb+YT4d5qkgNoHXqo3D8POYN/jVjeocPmZ3qK
XMzcv57Th2tYoeCRiVclyN6Z6MVpJK20hNAmn6ifxMk33JCYLq2ECZeHoUNUYKdWkOq8udr+JPF5
5J4lrSNKynCY161OwQETs04WHjSPhUE/q21/n5djbBwvS8QT5Ff8PVyKjUEvrsxPEhVvIxNTxISJ
TOT0a2/Uqf+3XQnTig1mshEh2XzMgeL9B+gUVRPNTGwLQhr0GWQNNbL15vDVrM/FHVbj3ZYSIohP
bVR4HK8B7Rx4s0L0VbF3hd2o3vjfEz8neUhvm/K9VgqNRZpu3zHqsM3TO6R9Y0CjZY7Oebpo4ZyS
7jnlwlxESSj6IM+RgYPU+xiRkSG2qQbzDPmyjTN8f9tVHZxvvMplSTlWYnYI8Qh2mHA/f8672Iu6
aPRaxQ7AoSDQ6JUxOyBWdfdxGmSxDlE6Qubr7SUpiCP69fb3w2PpegtDdV63u/u0gMjj6MNtL0iy
jF75H8LYeai/XkGyyaCPS4rdI7WV58AESImwCkdXjJLgggQJLEgt8QvA1hTi+kW2yC0KropRuYXV
BCEZtfxQ8MSi3S6/JLyWCmuNA001YHueSQbBLcTHxhbfa6GhH+zOQMmV2w7JTOkGUNCOF3MK6LKS
R5z5kbejYJrVqRuJHsmV6QUKJpOiEH31VrqhhHjeuIQpoSHczsSO5v6ijPIWA9+WycJ/arrwEJiq
wWALNlUT2pcWZT5jY27m2AmUuhZXJh8dQBrduImw9mpX07jhv0WeHBqdSCpuKCyFDqSCazy2Ijcg
1OBdFZZneYcJl74RHzHqO80s+Ad+ef11aTK8kfcSxtkIJW/9xXfSwdQAEZtamB/JAPkQuo42VgFy
LwINPuMfLF9cm756dsa+t5YhuXh4AZQACZ7ED0D97D+YE4zd3+lFhEQ1VZQTInehyYVZa3wUFy1D
OF/3me+f/WOaj1DdUXiIndxJY6EOpbIta/tx+IL+o0Qttb7zmUuXkbRPnws6FF81Ff7YJQJnZ8PH
cqhIqW9rWSChMGh2c6wqkaomb4sbDtr46Jr3kSxwsyao5/3VHV2KqUFGxHHsvuG7kCI/KprvBWCJ
mHjNZBVhp5n9EK3k1zYMCZgdO9+LukuD52aivLaEPK+kM2EX8OJmtTNYGAINZ+SbDtqQy5djO+Ls
SYkffQ0JRU3Sz3SQ7fEwGEaYwijGgj9pvn30BcABkZ2jv6fQEjIzUYZUP7kKp195fzGC46Z3kAZV
v0x1uGRPQ0TFHLpSaad3wCraUTf0zFLEKoKjZXjPJsbXEACJFMj7SJDmWpKJH+/EvKCAHACdC/Fl
A8KkaIQc82O1ej2kTYyFCyCXwH/199XtA3bBiY9cvUABMPWVvXnrZVDtbCcDAqcOsKp61fpZrLO6
MSeAA3x4je9cy50gR0IwtZR89jfvtY94eXD1DPqPfqFxcoqDIk3lIUtto/H5czA2bFETc9Wpm+Rg
QGVvUs+AqPdLf9greWldHmFoV/rcko+Boy6ABkdUOvFnrfxvB/CSv7R92KxWK22tIAjZG6DOLfHO
60vA1hLtt+5QoifM1jVOocQ4hizGlVqMiiguPphTXdKXbr02ikc/kzJFF6FI1IiMLPnAa/WSvI37
0K1ujexJzoTlUoMS8OuBxGiqW6dQQUsKEGe2dlY4vMmyASbcyRdHA31FxciHdyJ/W26NWRcgcCRw
XIbBkSdcV1clNGMZzIu40aVcAp47bvjI6fz6Xn7uDF+0scbL4OlaZzbtBsTOTLqgZIYfEoBolBhb
2Ov10oabBtQ6SvPOgfzW6AuiF8PDpvVjYcHovABUg7lxpH98kvLRFQaDicwOQsIRDeazAVmf0c+u
/zf/V/b8fg5naltZdkpZva45mEZi9EQm40mvCkOEn4MgLRytt5mCMfUzS4eMsu4aumhNTaOC2l5w
vY9Qsq3BsLVyVL0aBj2S4kTcba7pBeo6cssdlsjoGMbZr0ufQ7hLdN8W07ko4GQrhnHlWQo1Zl/T
Fl74BS/ypH6H0w5J1c0e9lA9svSETSFpUQzLYJncBE2mMLgtuf9wE9WH8e5ItumXnz8MpH30rQeM
oe0+YKnzWD0Np6XQopHZfJ3GbGQiiqNwJ8J5lXq6C4ZXqIkt8KUnmAjoIeu48kC3RwjfPYvFoRZY
7H2PsmyX2j6Q48ls5H06RqsHit4CeXuqX+12wFgFux9un/ItvGYknUhLOFftsCGDjHGHID3H17Ou
6Td/AtP1comGPotCMUtLvEjwHvt+fezPM2FFHULKaprGNjGXIkiaGAC6qhNLE6/zT8klEEzrte9I
HYIWBYu39QFvrAO8iZ4eoDGSyBE0NdyHq+R/I3h0gk1AQQCevAH1zK+bK4jDybONL+zpQD56EZac
wd434wujRWPQyABATSJDYuS6a/sKhBrX7qnRKPZoLv2J6sNWzzbANh1l4NquVG5LFuWrhc8L+lrm
X76FdFDtcqfig2/fDIuN/MnIjcCkQSvywbNkvfdxE9UTttPAyx2Pb1UW2QONynGxaJ6lvja1dFwz
l0JTyuv+JXKakgEJFSY9atcFjOAIdlZuGmk8ne1ObFCPSkxgAGK1Rizt9f9qZqS08aiZ42cqo9nW
OX88jDyRo4wuJEjQtfXfvRbREiFNZNF2K7I4HVfSfoRcJlIhGQ8hGXjxcDSJNZTR4rIyLAuoJ9yp
A5KhSCZAitvB5D0gH3yfrgjPh7JenqUWfVelBlV0pV/EmKs8HclJSsPVXJqCinkyC0iq37eUOv8U
TpvUoL6qmlTE7MyHr+CpD+bHSytIr0UnG0Yjy3+HVDVEtfm4BwyQAsLNMMrlve6MYCY/yChPwYmq
VulEsj4P19xWNbTcu3pIgv8YbbCcARJVcDw7q3XuexIhhFAGcCJlN3Zh0XCeHirJNHy7wGX91dtS
fSsM8c/w/6pRGSPO8WlEO1YMufOLgY1I0oN9CJzznurCXgxspravtfPYAc7XdKrZIR5UYTYQcMYH
RZXXXT8U1Mac6PyVr+hVMZEKb29hGGzjCcyrWQ28wH/V/RrbtTrtY3xeuXW+NvGMOZebJjKbmO4B
peEyM0hBoD0G8JbHLCXxDBsPdwDFjEGIs0CtXZsNe5j1bUUoecZ8lx1W3e0GgzOd2Fxq/T7zWH36
Ry1QW+C5hasNMGLRybUtCIPiAKci8UgnSw7L5xqLGnOG1s0oPwUE4Elzj/KiiRAtpz2ftitmuCyf
xOuviypLbPPYAHKYW5/8bP+srdixFmhxdnivKGGDpF4mA6VS7CksELSX3YRFLjLrA7gQ4i2gQAdp
XuVI2u3PKwlcYHAmGG7/opucuqhFF1hU9Tg0l4WgnrV39uP9eFr1hhOR82r60ycw7/tsey8r+oQn
6xvGrzaF4YG4uevesE4CNQBwM4nFfli/HhXsOyRqpliBNfCaG5o98y8n4zxKIJA/3Af2hnr18jA3
rvHipmkO1bCT3PNOAV2pQxsnqVJQOs4+z1+kEBn5qMukAVXTlUHhE5WXcFeG7rXPJMwmBQH0DQq7
RD7t7w4t4Kl6V5Tp0p1Id+vA9c5Ti0kDBAL5fb0dkDCzveXUDLaqi+mDILRheATuw7MEgCX92l6B
erNfqbf+U8XLIG5p49/yAi405ajd4eZcHTxpF3sbEGAL/iltqEaqqVGgOZx1D5hWjNYHPn8Xc9w8
9760fBSmgtFgv3jvUTWq6a9d7wCY+t8bYFuD/XS5PIr9FXX1DNmVEHjxnreqK1sw4oHBK4+/sJh/
B2BOe+cRGmfjrkLQniZkDdnP+gsXAdXgYFMmZwNetLBYY3X0uGLkSJMrcq99KGfv1n9mbnx1hNNk
cTAdM5xGLTFbXNRUD2GWX6cq49J+UpWti1rmszoqttGa9gTdnfK2IbMUL8KTzCVNvIiTxmxB9UK2
UmNx+GrwEElQxC3eBtnydMyjpBMLmXq1Qd7bo59X1xMdJAiWZv4DuZte4Pn/GCvJ0ONW8ieZQbJ9
IxkROljleAd5nW9LGwd0jb0sfUzUkVvmlW76X29K+33UyimJpNHFOlGASwmhaIB82DQg6yXmNYg8
tQccykzKleaSWgLMFY48V55h4Ozu+lHBnl/J1y/DKlScoEFQalxj//yCex/I3ypkr1h5UfbqCQTz
yt2fAjucwrfjV8yJjZs4O9Gi49nNHBVHH7moTec0+NNyeyJ+xSTF/aAJKh/jqY7a0Jnz2F22Q5TV
jgDnvlHXde9rNY4fogwIZ0jfc8fcYEkGAOGP8daBRP9acb+5EfTexvUUY/oR83v8d2pn77NeHNi+
Prk734DhHbOrGp2RRHo3ObxeJChsIJXtTgdDLiNJ0Bty+/W7XFBEeGpGLY8f2rwXPuyX5JMV0FL3
Zv7rbNOUh9OA1CIqTSpGXbirzTq2D7H51QqvopiOZxrp3aMRl/pkF2Zqg6jgLVRoqNtBiwlNnH8f
WRxC+R9v2fpTo/fcTjxE2xEuiunWZtF/3W1wNNvafgcwrQlrijC12SISf4nTeyNj8PlQqjcVohTv
6LAWR98Lmv0UXOuShzXIVSrBDOy604EI9QPPClHbnMTF0WwxllJUodW8BCmoZLpe0k6asDglEthf
gMliphV/JbjIQvMhr0rKAuAtaYbSfa6IoK2XHlS338etSHe0QmboeAhLIUBTmE21aVpWtbXRAQ/G
GsE7jYSwQFYcUnMp73xQetWS2e1ZxBv+owDLrYih1Hl0PvlQjOacQezSYKRgV9AwzsCIghpvoWrV
5+wenXLG0ZnhlbEY2pwxT09549QYbB4FrycfVkG0TLo4B3GBe9JNwDPp9ikEXf/ouyh1vLjJLs3b
kwuYfFPE1Uac4QXmdw4bgGCo+d+rBScQZnhVOMqpG+O3n5pukq66o36wZa/bjz6mQGUvIs8ZFXlq
5n5i8+8sptz/AG41/VmIUB2NM7d7kPsYhWnJy/cXoBtsGweSvZ32U7mtBo0sm1GzHPBIOlpJgOAr
wIPYpRym7u+V8Q/fd65VdLgyoKVSSmaYvyeaAOVpq8I4Ddb70wjLhodBsUUbX5JpNT/HhYayiTOp
H0C1tiuGRHdxFRhWSARVKk620Ugds8lz06Gq+cpwGUfXKET/6mE+NGlYRH8ectk+aZ4jqlSoD/sN
PJqlbPz53PS7UgqgsAjhvkpOQG3KPnwZnX8Koh9i45YHy6DDGIV7NY+FnMdtA0GijVHixTYtbDKN
Sen7RxCMg/NoGkeKQ847OROWo9E4SckJw2F2MqUalpmdt63J14kMId6JvATDHBxmqwFHLm99mWg3
yV6yvssDz/J6cgcE4Ia3QLAi6CPKCucK2ulgcX1BrNi8Et51f3Um3TpbDLT0o2PLrvpKWlWYCMfB
o2TeEtoe5/hA9Nho4o1es0NNhbByxUjHzbnq98Rey7uLsb0lQVDJdz09GjGGRV+j0GTD0FyDRlui
EHOrODmrcODqwFPzZP8jRgyJlKhNgFoxkgz9smxu6T5BO/ytzjJJ15enjNirNDEYGrlTe5uRS64r
SCnI4bN0d8WU0N5RbUxtrtM+AfDTBgwdU3V5A7kZ1SJq9V2YjZv524mm05ztW4eQ0E6/dlCE9i28
jk0Ediq0B2wffNg2fnYC92dEzWDIPsspM5du+tHIKRGRb2k0/2OT/GukEIjk7eqNZSfhWgVAy3Zv
4Hsl3tc+62gpvHpbiGyaPEhXcPujrz7C//eaFsPKb+1Cju3k2XLEKxSYmPY3uhtgTs3TzUqMk0xi
6LJda8b/jzWhXViAZ3qiOriwxxK5hCh8WBaDUwRAY4N5ySa603JH9oml56cPz/VwBi/KhVigz+Hb
ItaW+FMiDmd+pTjaeyxgvLOf/wdYSBDJMfCYtijWC0GgF/0eeEu0TxA6Yk3txOxM+jELrPXvh6oW
Mbl4ce8tWNn5wtfeNosahDiEr9mtMjOxGI1N3Vzuh74CpTFJMipkdAUHxE78NtREvoTLzyOug617
nSM91nqeUrh4PW6p6uRlHZQQeB2OrktZ1efby1TTWxJJOH+VvytAaIpAyWXfCRWoHEIW/xQAK0uF
fHos4nceIrHFo0wmnUkIJGDmPOWI7gFnTFhOiRYJX8lt6XYx0Zo9Fj1IP8NzDKwy5r7ITB07q8eA
OnNq6VDF4v0KdT69gmfmcKfM4yXx7prr/H6gNlQDc84ggwLM0ggkPdH9TIgdxgVGeVmb+kIkoAXs
1fNDkpCbJ6AbejZgaq075FeMaEvdvtt+4o5/aBUUXBlbmHBBBI5L37pTM0Jm4LqNZUSH6LrRV3TT
W4tJRTGNbKDDgQzjSyDLW1l92TtaJdqBBGQaVkCDJc5QZsLAKZAJmCE0vY0/Q9RIl8mp+h0fQt6r
3ahjoY3WIW4+yMFvyQa2AqyKZJkJ+qWDevW9g5+CI0bJFA5MviZB3IN0qECUSiLdjA3XBCZ3zaGP
I2y9yPyBYENtvaqVZVlkhGoQQzQ6Oe/0WWbnMOoaNHGdLm9HOKta4Nc+cEvQsf6UtvR7wDjsgJRe
mfx26hHp9VB3eFCAul5oKXx+THYSd7j2dAfxaJUQnpJggE5wmL3ArHeAnstbAouMMGFt+633w7oq
Dk6iOzCcDwKbbDV6YtTOgk++xhmJVb8xvF/CpLPKpuB5CW6f4z7mt9tHbgru5ZXZKFVY5ko+VpCC
IDY5/RiJlt6uG1+xPggS+6WK13MkpFoWyFVKatXm2B9P+b+lzRrJlmWZvU5HCSfMA+gnPLjS/M9D
fR2Tr5poSdbshrE+mldc3AenDyvfvwXtdlVPM5Kk6twIHIbuaQDNbgp+Xuq3Om5Pb33QZokeSL0J
8OhbPbHjhTRxZNNqb/l1EGiY27YnbpdXj21DNnGrypND0ONu7z/GG9epBjeBlv7ql4NQvXZ48ML3
fZQDXgTz6VrW6Gswt+wecYvJrRUsFiX5/3iQ+dJJWUU2d8EOm3PLzgGF3lMlgj9v/+xRPFpO/+p5
6iS6Sj1n2rzh5DPpnONeR+pQkSYhB0H5aaoBdPajJPKcV5ZdM6Hlj91tnsBHKt7w7QZ81VtovJ66
JddlJVdfR+2hi3y/yc5otAHBnVElKvwQNhCNLK8hErGLZnsA5CTOS6mD6gWcr5vo8KVRRhp4Z24X
q/Cqfmr+Y0xDB3RA4KnsXHWjaLTmug6wewbH2vJr+FIfETidaBndJcqohakoEZESWmtCwcPydX5n
LzxNZjU8f5TchSHO3zu7BngdWmw7Qyutcr2VxbK24DszP8lOZ33fsmki8bb3iLL3sGJAzMff14bG
QmysXaMt9WJIyWv9w06xdx3OB2cTklndp4dWPVveVFrrX0DrocNBKw6E8WwmPr8PBYB5HEUCxnEV
0tSrX3bd/u/Y+OCyYU+ROhPtMbfAY+Y8unhFhqt/HGnlzDHKJOC0PjUCGnSS2Rpb+6bowURA3Stw
YxY/B/ifqEgG48MuGz8zS1FCsHb1Rj47coIfZ2n0ZRVallzl/Kh+DIh6PxYLMgYAgdo/dTDWRGib
70Blkr5GkeEJAn5bWYuGmQWgi883sTXTbCQjA0JOvYIrPTOYYiTfFAIdogKGswQ8WWMfxGnbTjXE
3IiofmDIM8OnDK2lIxm820zb+kCzSbosnSl2pHTmlExZA/3KMkVnAm3NL3TTIL9h/3iV+2Kpxr9O
0xKrYFrcbs7ayQsbaBhZxvv9R5VjC29RBad25/Y6hx0CGrFjNvwG3ic2dK1PNxACUL9zZTljNoKq
RGq0ug8963+YvaGfXmAINKKWNE21pt38XJdtXzRd9faYy7z98k6MRmck97a3LZ8WauevrZ1CsqxD
tZZw9QIzPrBz7JGDekgPo/jJaV9qXgU60AKSvLXx5giDYXFF532NrEnu6oS9/9cw1psiheD6yz/F
3K4yZ3vPIKL2pCPtyGlueuHrihMVI29H3cEM14au4RE6WpWgWK8uDxBq8PDthIGOWatGlvVYnUsY
QaPjwKYefMepsKjWdYwGOGGUL+Xpcm/OcuRrTHwqwCEQdNWU17gjlHLu37eMXg273OMeE6zddr5t
TwDA5maR7tJP5/KEFqgColN1jiz2LFqCxg1ftLH0ix7yq2plw17vvpZnZM+fzlI8WFIVE9zGPHQ8
ptzHWR8P/t6+VP1itrTLdb/UK5ktRfo14VMG2mpMXdlIX3hVdndhhvKKkHrT/J94Tb1QAKjSNmId
rCgqaPabhiG4P0ns39lN0469DJR+k4YnRpRPlnLdeakH2lTVxDjwadYcgm6HyXu/ypJyScnVKcQo
S+ELnkSeAlOsALE9OwlmnyXC0uTxhspg6N8tFjMSm2gMjma4XKmB3u4UYmvZ/dJIEL+qcbTJBfp7
yBNxNJXwOGyj6PF65YwmAxdNmzMepGiLVRKjqrPinAx3W8b745WijNp/VbjDLIsOtS0G6cTjxdRm
sofWzbzXtT3YitrRLtgR/cmBSIIKsNSRsQApXtgE+QO1/jv8VZQWgmaKf1VGC5OFg8Yyq9qetfQR
0mjcPLdaBRJ9Pzam4okwX1b/X1Ca2tnZORQx6Ql+fZkDkxrOeENmRMw0oIxSJ/tksvttJooa6sp4
J8IgaC5vVi6n8hjq9ClI5lmfOYiIuaRFGgXdmVMT7w4fi3cG3Fb/tKZtbU06xvs7wOCLF/Y+F7MU
DFSZofyoV2u/3KJC/jiGpEZ3zLz5+fMHkpNs6sMWxNrWpwaQUyImRpCVLuHII9EVpwfjJCLg/uVU
sP126IoEf1R2eTEw56f6yIcXe1m6ZRPZtDVrqNmkPshWV3llbZUDCPop2c/PSi8/kkW0+zq52WRT
qS0wM/kVwLna5P3lMwH76BohFXaj574avrg5NGxU5IC9laqGVo39W+eSsXA+c7NkEhOoah7oX/xN
nSYDYoWO+YXFlGclD9hSwkabboDlnMknwx/jU99B0Sea4WuBWAfWUqOSPWzRH7jNS8SFM4DfV3aU
wKxgu6Ez0SeCYkNHWk0AkOiX7Kw4SGbIv2wdMqmWh99cWb+McTJtDc1AJLvpPE97dgBujeO1K7LF
wtQ5oBK9NZ8aXDjWxB/UxBhacGvBV1jZcPYAwsNZm7NDALOSvHGLjoNO1CoFXdutANagsa7e5Zrd
LhE9HOlp/x4kkQkhnMAyjYoJce+cY6PoHnG2BH1w5X+X2xGBPJFhzcxirDGtmNHxznQ2RXTueHM9
pUZMqtnqnGacOmv/vwpc0H/Uohx2DkOOSfwArcJWzcopiLHpxjIYadyBHVYtWzgDS3SmybChEqNC
99GCediH7REGCNSHWDMgdDvxxdZycIEvdJR4idcwEZXwrZlHwV4FgaCcsSXuzNXS7eSutRMr/nns
EIFk+ktoZjV3CD63Qr1Z5jLGP3w0QHYrXwxz01ymakYDYqr1/n2yvJJc9rlxsrcttMaPqIyPanqg
sUsfMBGw+JtFJUVs5726p6i2Yzzwb9bzBX5M+QiYMaqCd3ZF6VnHioyxB1BBA03a4qRGC/ccAGUi
xykPiovgsWIiUjxQOViDdEFpm/Mcw9omDFkB92YFvaZwrK/wioH4iliImZ8+L7vDtnK1QbUUwBFD
XmMrwfMtPW0P0Y39vgsjgUcWEPt0letS1sjada5edtmbb2SBJiaseBgqVFPfYlQ2ZN7ZcfU+zwb2
3WQADTfN72O3hzG5NozfXVgn7TCynOi0ynVGB4zfIKXrM/56OjKvvHyrX4gizOYKVXbN6ffl9IQW
r25Uj0sa2YvIKiWCjy93yi7qTZHsu2EWqfsAmofe4eE6RWTicxPFlFybsLsIJcnvvF3u8nFvPrIH
EYgltD8mKWDNL1gGEH2zIIh6jg75x50QOnA04mBvdbTDR8Qv88CEofeIxGa1xDUOmv2Ta+zIGEax
V0r7FM+Lg47xqn9pup/iCR+uykOlngJBAJ4IEsxhWkpjX6Ns0HdthtSfderalioE7IX+dQ8/5n7H
2VyvV2MD4v4C5myCIRa+icqN1rHd6VrodUr190n2jiL9XwZN6sWXQYD4EFQJglyPixjKfh3RW7cI
EKKJJgPTPSzpwhVqzbC6zcRwAPg93Hq0+NMFDmD3xtJcni3slxYIwQUTKCdUQYei5mVgXJdlHQ0D
bSVH510yWSoybyNanxOX9vjVRxse4XsLPMXQBOWyziN2/dvmbZB7fBB6z9BdakYWF9PRW93DHJRW
gSplQ9pVMytCuBmvbT1niRc7fcprRwTcUltIToI7zO0YvuIC4r025Tm+99kchsTeK6GjpPU9nJIL
kegbip5hbXdhsdmANHzQ1q2Bww3nYqoFnAH5aUh30/98nA9osMUBwJgfDfwvsekh1B9CtfqQxY44
l+MnGjGkrkGU8ZQpPYMTHIesmovmTtOlGk4xmPAjtndbojEzMU/Hw2yKCSTaM4DjECU2TJ6tW+Zi
AnqK0OYREuMQ7LOVLiIWHZ+69a02C/zKvvTR+NlvfUFvUC4b9FOuLZDvbvMqbXwLNJgOwi1MZMmB
E/MfjDGPSom2Yl5qeGMCPRDwYoK4gk/OKpAhJX+NXmQjRgE7d8SCS3vWRgTKFVmZdcUKt3XJWH7k
yXbjD1gyZBsWyMzH3WGoW56lStaoXSbo0z6Qo1eDlnJhKfrRRpibApOSVvb8rQocZ+OQGU93iP3H
r4/bL1GyWyYuUPjHOC+82GiGxVWtDmSktLIVa/krp4lvgsV2JA+BAxQY3tRQxckNJRA2TgGRPe/H
2+cRXoEOGP252Bl5gAeNIkwHa2mhqxwrdRUZr9RuJZkd5gnTBxPYZ/c+ghPaJJsyOK0xgqM82GGs
A4yIhJFNykrAObDJk3rbICCCF6O9F4UnVxLlDWdtUpS2JUsByZtdeFpnRHxonf9pnkx9RKkolu7w
1UEKHULimDbiE0JC6Gva2cMY2Qjf8VaSXTqNblVGTdCI9pxnvbgXr6PiDnnadJj8fmQks4oQZfVq
uxOSJ3IgK+fwOMrMqqIXRxz/kay2RSdiBUSyop72s+upMyQWQ6FdOQSdv1vC7vYpliJOVoXBKh0l
BQQeBMGikUdTXfXA28WAR5SqMWW/EegrQigVTM08M5Rob1h4QwAA7JFWKriU9x8HJpANRhPn/4DC
rn6Z65B3aOhWE8mPsQgFvPF/JRP77OLZ1mvQkcx++6HBVB80n5yhaftYcR7uJM+yuB732VVWUjha
GuHweEokZ5EUbf5EMrKTXrr3ZMnujzX2h/0b0nlXCjDm/pC02BqPkY9CjVIVJN/WZRtWki8Nir57
W1VjvGr8ob3Ur7P6XX+GVsR53Rby98RLs0J8E1HE/Teshem+y4CZo2RPJuGQF1YZ6SNuaE8qqUy0
/hCrizK0rn1EDIPrgGFvdGVqgGNnD/JNQmd5Al7S0AeqmYFk9HgAKrufpy1x8P8ZUjnD0I+xnJqc
nojNFvucd81Sw5YwhaYXqw4ZkrJmwyIU97A4PXNrkAu3EJe5KIkhDBI08yggbH/YifeB0gtiXFw+
a0vs/t77f0wvsm02viFCDfe4XN5TOMKuhBKl0+eZ9TzNtZBAodMPp47Onh7J41rMeq6kwJ/qSMUN
BrUacs6JFS+dubHKYss8gznQODIyxyKsuHdWM8uncWuYak54W8zu6CPRB7UtQMgc2Sxe5GxFk0aF
++1AaXYKzH980YltKDglLQEmBv5OeiHq7Bxv7EQDxfSbRfzBb2yGqpYiIrcWnZkILbjvOjidQku1
X7G7knaKoazNpIdypz48kjCvJUTlESCdY2XSgZTZE4yS1NYzd7VlPpA9pdm3y+MrSUGMJAduXbeh
amCw28h7GdG4EswkMkspv6GLXW09NP66CpUf1vbiwOkN/wkoDuFsKT64GvSHwrt2tewmMMXoGi8s
dzazk/Om2XmwU1Z9h2p+U/Nt9HJzKdA5hWbPwdiZOOuCmZ1tf39fNoheVAKLg/c9RLbDDq306RQv
kFI3rGd6YHrzuDwMMvk3NEZW6+zGu/5eqs04dP3tyy0wHJMjhDEgd7Syz2vt2vqlGVsfyTjQH0+l
KEKDjYG6SJ0HZx9qSk5Q7dRu8XVogVIOOOcS3IdNuKcHv8pqqlDVCGRLyOtOkoLWsOBAJLphF/2g
SCNJOnatVhgL0OzYHcYwluQPzrnKXIKXlFodpxd8gbL1fLWlwklB1ox1wc65PTqOl+YfnlrTSKW0
mQ7/gfs2xP9ZMnr4P2bjQztRkjtfE0m2mmxzQzZjcZuNNsE8lLrlCPreQp3lNHhXA3QfUKu5hfd9
QQJE3RtyvyPNoDbAGQc2vCR2RpUpTadzytzc6daau0lmnx7G1wQ008HYhD+lMuCD8jGmamG5826C
qiNgV6AEoKD3TWgYBlWrb4YoDY0UjGMcX3HHes9m11g0WqcV3zC0JWmpi1VDZIA6vnqZXfunsmPu
YSy3LTqtV4FqUNAITGFkVgp1gtPp5y/tscqCidXDAxaghQ5XoduLg91Re8T4Xt0NpzYkWdOyAmqS
zVIqzz6JV6pXat/8j4IUMr8ZTFuZx/R+sK/5sTvbT9T5Y4JwZ1KLZ5nPiVKYNSufEhzFdZXqfkho
YD3ZPKS3twq8/vr64UMk+/nKiKURTx40BDdzI4fpKiCmNMR3nqSXoPN2DjS66c16THWE/Q5sPK/t
EKHU/L6NEHvuaebDc2dX/mswNYb1wKBUUq6sI4vhoXIbdjDPh5D7Cf/I9rHI8sjTSj4F8TBGL081
JxVQhvowspteHRMHRv4S9FQUVdrcjAtOnMgaVQg0j1aXTPfy/coxqqqhoqqs1miS3oQyIPnNPb/O
YrRnD7msOX2aBy7U9BRtd4vA3RE73gNfbuVMuXqmTEns5Hc7snzctGBlIg/Nu3OLp4ks+CkWy4o5
OolNXG8IEz40Efr/vGndM3OIdavOrUdgwz5ksafapykBGQ6262CWWCnZ5sH/aBf3E0fTGNkuHUZK
ljjytuJTl+aqS4hTtghjqM+IG6Bjexhg7BLNSsDXULFIO4vm1vSOOMXGaqKoZ8f0kbhD+DsrImmv
P9n7GYbBT/gtqK82pTHoNlIPSTiwSNmtxUvc4CfBqkm4VoLttv4WcuvD0sapA/on1KZYkEzaZV6D
kmMk/HDiQgOwSHPtlcH+nlAVXi9yz4HrU8c0xMnzEepkUeIRK/dN1Kt1tSkVuN4ds2b6TCZ7/qOi
Yr1Fa+mpyLzB6ept6uYs7TinruKxFNFdtYpY89UIFHxXS/HEQ98Ke62DOHzXP0o9qnZc2nR9jyA1
NSv4O8YrUwo+gY/Jq9tjARln6QNo62xU2uSTTPBQDPy4MHQHmwH2kz4ScBD3wvv39xEw+EJkKRDP
CrjBs2ZoZqww7vWJTIGZnBnnrlyk1/18eS9gWFkkpTsuH7vENWHR+/p+877eHW7v+cZ039YXh3qQ
m2d5poRIi5beEGxLLcCwQ7NnnDuFSM2iXZSuoIL5Bm6tMr84bBfEJEfIaM1ng2W3Y/3GYFaMPDUC
Nd+5ABQX2WRxx9X61XSuNnR9b5t6pv/7+RV/32x+LzCQNoaQokh3rl9wvlwMU8sUYp79pO0b46hk
Fpnmsombvs8jTD1JZdn7u7AL8SLBG/5bKDe4V6b4aoD5TL89+rtQHYBfDhup7At59PWZceH1X5vF
c9nmdkIaVSqLCKopV0KowHNA6YvA6tx0D8gsKi8hWH13CRzJoj3vmJNL1p5SC8MiWHZgN7eEUvvN
GfVjzD9tqf7Yw5rUUVO2egNQkViyZdAX3yeOBjDZy5AoJ5FoP+K6AIywyrEjNTMX+dzF+q2oL0mR
mGLpMXjIKTyiExfRaVGYwr7y7m+yRmokhBve6IrckKW4t0I6evazjdNarWGuXqsZf6HDfwN2AU8m
gmyTN1wF9bn3rKJc7OG/IY+mkXg1SEVBfkU84ptRkox4WkL1Wgfg29WifTUYxCVQ/fb+E0QKiiba
SEReDs4N/dZqSFmudSe10Xk3rJ2mKh+856Q4IvBg5NXgF6VwWQNW+bEL07H1MHnAs97ErVG1ruXQ
rMfPX0obggLksycl+DPYh83MeDbMdLC1dWD7ukuMe1UEj7kJj3R2jOe6hvQnBJEKvfVT7E6S/Q2f
aYDgXsHrFVPE+fFb0YqLlNJccuZV5zHWGwGMS1K9AKOrI/rxx0YZ4CvaWfWriUguA6sOXtjbm4Dd
BZf2RBkngw5vir2ioE6Gt1yWjJJV1vswsHP4cSQFQVeT0sK1JhbAMSK9CrLFVkdwteIsueU7ATzt
XpRDwnCtS5VhMjMD6CdsEolRZzaUmyq9mLsmW94Tqlt6iXZS88dduM7MYJT+SK6mweZx4rs48WDd
zPbr6w3RPEQeW7ocRaB3XkyEPfgKFCpkB4wO2dmSEz+vozOu4eSmyEiNqX0bZqbDGk9yFIQu8dZX
GwJ8iPeYJ8S0r0e3sbAzc/cnwhVxm9b8riLQm+y6xW+2enyXp9RxqVdwO/IzFIMHxtPEnTIF7ylD
KjQ0Mkvot1y6dbxxIpNLVgwSQYBlVcMjV+FiG+K+ardebtthUds0qRiAS4mEfeP1FWDgk1NiugQE
InBF+BEQGYXe6AnX+pETXc2C+5NJgGf6KP4pRcXrAhUh4owE5bc8vw3z+AmxmIVTNklx/MoIS7xW
B76lI+ET/fOadx9saaBqcxTDvkl3UWdZ/MQIC0I552Bd/gjN0Tev85VmNOFtsFfLhf2jFxFL+A0q
95lIPTG0LGOJxDF/kn9cAcqU2w0dC/DJY586TZ8jYEq5W8j0cMogn7Zjit8XagfHAL4RPguldEvR
q7CIBF5Q5dYr0XIMa+LsvG70wca6yRubJDKTYHWvX20/5uDXGbWRrN/7KQMzWyfdEdoM7fOwFMau
xhL4JHvOywaBtd15FqNtZR1HPXS54RSfs+R/ncQJgI/7EG4Qrw6BialtmmpY5HlPa6UM6smbwj/8
ipEU2MXUOWRqqR225p3RyVEMN/NY1dAf1sGNpJX7fyWV9BGsvfi/OxJIw+JcddNwnqPm/9OUmT22
tWPij8CiSScWLv/SHCJBCd+2x/fLlyw9Bd8Wt4O4PJkXdKnWAmVn3lhuVxCPKwRmqbRE27B+QHgZ
pIoznEuD11zewppbkkK2CXt2xr2CnB4K9hNANBqFIK4m1MLAVeCuaa0VbwOCobHoZREVxA2nW9+z
TKJ2Rqa0/pCUoc4C8xEyvTdEpvt2bRykytfrbtkimPVEbKS6bME+SnKIa1mG10ekWsPedcJI/js8
FvU+ZMY+JKLPwAG3S2lMWbRUIiGH3TEZX0RqqMhe5C/pZArGNRlHSy9fUzA4/g0Vmoytu6rivh44
OqqTpB0kFK4ecqqi0A23sF/zfoa4iTOHXqom2ilOJCBX593gCaNPwCB7s2EFMVkN9ukd+Rmx7GpO
zfIXve1NgsaO2y6QAfu/H94Eghy8FnjlKTt8DGrWytTj7jqxAiqMwri8IuG1YkCetwdb5dBQdrYi
Su7Hu1QJ7GkEXt549NFCry4WtdGsBRtatzutNHFuT+o0W4uHfKCjGjYX2joAovu7pFYdVMo1KJce
xjPqpDrRCaKWT3P0Cy2NaOmSNBZqh0A+7iliNAQHZohG4UAeeEy2eYsFWr/LxyfaJflSyFi8WyG3
Ud1lKyOMPhJSlAbU/9GzGlrPkma/Al4GJlIciXi+7iHvrXlfZP6KpPuE56GMmReUKJovK/nN+ahw
TLcc15hBzq3huT+3o71sq+l2P6jnho7XLbZRNSlADKA1iN8ujk62Gnfoe8HKj/FTwYKyQbHQMNiC
L2SOwyiH+WJdvsQCbT8Vi1bzPPGmN+TJgCs6Vq8xiTQSHilSbKcAQOj5Ii5OkEdVQ88FsqpF9IYM
HomUY/OsSzzUfEsF9k0ITUgsIt9iT66qcPxme6TmGDKbDURDXMuUvdDxo5Cc/i8u1Zmka5ft9L4d
hXZh67AqujfM9pvgRLe/8HW5ozA2DWywdAlx4BaNpn4sBHzONvbcfzJWUMvh1nQZhgzimIDnhoEw
FQyuUmUphHwHOFqQnZNoaHODUDr2KT7LVIkxsL4ZL5yR0HGp7Aj0tEBvT0+9oPX8E4BYJHoHe21k
cAHrClcl4mOjRCK+fQycZqUv1ZWOWu6EQoIDqsox6Wmjc1gRK7dDl8wI4UdgXzVCrT4ZcMe2R8iS
5+aOa2jYuf9ck3YsLQSnhoSTN7D0sTg+CoxuB4xX/DQGu5l2xKrZlJrz3401smTYGKXUFPzqg5kv
7B49iINRI9gHF0AcKvdRmCTX2vki3zLiC3gAzyOfWhHfiar6ZWEXLXYZi3pKVzhmLlRNYB5CJwam
eLzRGfPbYgYokRh9cOufYR4Ly7IyjawZp8B4nGmnf59LqHTrCz3NqPkJgkMqLQ/+6dHqeKgSXXiC
03b+p4Odttfe2mfMhOz0bksa8w6q9Ja6PGwDL9O79ebbFMayGor6wdxlOQbNN2UzCmOOhbbAzttK
WD+3kiQ/QdCeQ2LVqG6+JUwxgBE6zeIEKvMPp8YbFrQTBBQfm6VlopiDdPQdm2H1O4mWtHB9OY4y
MUMv6Ejl9yvCFUOFWe4BHfxFSkN5dMyr3/6lcpQMtfNhnOnzvKUYAcH0tH2gIEvVsmKzGJjTQ0Y3
ARGzACDJa+YShFY8F8rYMSEskw1mFJ9Md88qh8E0DfHDPZF+QyY52WDepX1s9LyVFZ9jwVvYBlz8
Sg+uVcqA3w5Rs6kcOU/JDQ/US+RBKj1eygQAp6X6b9ROnhOxPxkh879j5xNiIeV5kOfWysaKeIZ9
/H2aHavmUp8Q18ruidgnrS2hVzE+eqoFxKvkqPp9YLF1EDsy+B59sqhf1GZKhOOFhCzpbgin/YoY
k0lehVe2z6rbrQhUx5WKyRRrWkHvqrRPHKKEp/U9X2lRhqqU2C4ySTa9fLI51r0V9lSbU6RInRnq
qEX7Fb1+ZGHPO1mFH5s3HTYV6GqgqlyyuU+MSD1NDgm3z0RrUMDpC+KpIl7i47FSUXrFxW4aZUaK
7VHt/mMM8QxJbKjoSSwEypaiBLwjxAQJ3mYONHDUQkelSRfED/50sP9X/IXTDh9bGJGbAzjHv7Jx
h3lxnFJg8iKXeEgGkXbmNY3fH5NAhw3jOCf0kWu41hwblJj58kV3d9dbkqZuBgCr+Lp5hhZU/NI1
NNh9jpZUdzQaA3izjBSDr1zBn9TeoxOvWQOWIRe21y8Q4guwbgDzG+CWHdzp3XEHs1N/+OClOdL6
dwkJhkURpkc/XkmzKi6ddajqev7hOlcwN5disk/emV4yl/3rweOw0N2RAaFu8Jbhz5DWKggXngNX
QYtOr/47t9WQV3r09R4ixAyQo0wsimJ1f+RF0bUR1njffJ1HxQPqKwHAlvOFL3rZ/91Tym1+/Ch4
CWZz9EXnRuSI7GD0oMkO7SUZBuq1dP60IgsqnoS4A7tmmsJtwQ4StpjLbxKDW6VFV08DULGh2NZ0
97cD9Xu/gZPrsyRp8GzGzbeEiYTzxffpbIBI3Ezh4KKIdw8B4ht5V8bKaMzBoSX9YELqFHk4GjGx
lj2osgWD22wNPileOP6RltHCKyNE1ZEDP6nLT5+Nv7+zu3DDRNDGym8EI/4qXhFszS72w6tClfFB
ZQNt8IqzHFOws3dumFX791hvs03glXrPBVgmgHzkQGABSuy/Sn+HKGfIJJePVd89FmRrkcZ0+fth
y0tzkajWIUQCOuQ68sLn/MDdOuX4BUXAdyfyUYcPY26ZjskN9lc0qdKnAwRuQ33Z/t8sIE28+D9A
c2oOah7pyDDjXaEMCQFCZ3cIGHVxDyjYE6oF1OfnnUT4GwcDxQGpJEnpxgwTmhNEiBcV3sSHOavS
r/FZPNYW7B7cyQBq5/sjugoPbXxWsIZXjNZT2ughaM2X62izmpJhsrxou1O+c4R3l4y4EFPXhhHr
59ySAKEM5TcSWzOAznjj5vlwgZNUrHfiGu+AKRdtPUGj9YaBgzuzGB7dq0SZGQHwKu3HFQBi11YQ
inTfONnk9n2BzD+Rz2uEcJYbScAHaQBf/ofpvYV+36ol5yhvi9f6Dfq8/oqv9TCRf7AxSyhR1Dwo
MCG5pE8K9oKYFSqXPKGqTiAXJ2uGtxk3zbDE6EbSnroAD1Fy6zPV9y/1QjaG4H5dNGGLkWV3EIja
uw/Np+w3Dkuf4W7ZBI+3YTof5wzJZ0ds0bScH3HHrsM1ctGeZUlnj/ait9XzEeWw1rJkD6UUD5V7
g8LPE2mNk9ZyMXyb5vj9vxECtL/6FJ62q/rAO/MKmeJzA7YQVMY2P7kpEUFe5OJDaf2cra6e1xge
dFxRV1943JTn7hJ7j0RQEDM3M5KhInwC1CfskSkPVBoMe9ds0f/yUNqPrBgb3n15J3+hASMlAWul
XFHTgRXcFADO4HkPk2VZqJs7dDNJDPYoxYD62/gBnnRLY8RBS1x13KSAbI2+t3VquuLZqndFDvP/
om3K7IjYvOfG9d0mgMeTmdfdAN5gebKbXvEe++GuE2qbULdnMHAFZsQcYGtgfMy8NBYstdpym/AS
Xr4JDVyn+BQ74mfJKDj+pACpg0EwML2yuhV9Wcga15F1Xtl20meZBWvaLEZY8CKQfpodcmHkq4bs
XNBj4v6iNd5DisfHAJBDm0HKP9D5er+FSrh73ZPIcm/Odm+tOEddqSWORaFpPyfqG2Su23C/QHRm
Gapu0hoAHRQbCiLq7l/rGjfgjR3u4kwm0dY2RKM6/1+OZNAqIam4XklUSehYti+ZfuCtCbDX4I/f
4TY6ErkvDcwgASgyvQUUAewGaiKl+HRecnZrDtzqqdjalVzznJtE4l8H9kDD4tpy6h0oC4+4+/+1
WC4UQH688DdlPgj7ELcDXgCA7Pyf2AplunHRSeCXFpO40tqARGKvslNa3//wh1JdypOlGsxxIJv8
lC9KvVP1VxGxq1a44kp0jMCAAsTUZ6q5Z3+M7UnLmVm/+FBMKXj5ntVIDF8OeP3MqGHxlagEPMJd
BrhLP3g717zhjo4k+ih/l7ETGpYOV77Iw7K+vzIm0yaZTiNtQqWeI6Ieox9qx813iitBj2KXn592
ZSCJXmIxOXkvROnRzCKNtFSbTAMcwOpz146hykeL30kb3SNplmZaxtPZn6V8enbizUg/QIn0RMsH
uckMvpdtqacRkOdNd3ST+F2q0hVOSXiIOtXjbz7xBJkq3QwiWF+C80z0F8pjEmehrNRcbQv3F+Ug
uCjlA+CraSV88W3ejd34PbBhRc6SW+idwRg/8fXax5czBD/Px30krb+apBb+4FW4BcFdaH1szKJr
q5fMrhFXvqWgpjam+el8CgkhFaIROowB0KQ6MaEtCyViZiQB55xRIjZ+vxYpL3SbT+V/INKW+kYp
cUUW7Gc8Psu0HLqObFuRVfEHbzJZeMccyBfwEwV2EQdIDl+Rs/7puUgVTdvG6PI6TK+uD5lW3PbT
d0odf/UKWVxQ6DQOjgJCBRFN/G4omVypkC78fRijtDSO2ssMHM14Lj29RugqT2dhzw63aYuyR5XB
Z0QMJPc7dXXx66X1ugkE+ip5xjDWTNmK5EOBC5fxSp3XIRYEinsLimhRMKNIC8KPkr+40Cog09+k
Ba4FKkkG5IoAmcdElwGkSp/j9wcEDP0nIvv6iwRFJ6MgbiYud9BahovdqYnaIUyQcx6VSe9a2xVa
jY+6yRBQ8+ykNSEL2rNg6ceUiqwrIKSEynyg0aQzslk+/V8T8k3e/R0vbUfjHhP39/jSp3s0mhsU
b+yItoZJ+C6LJbu91FLE+5FQ1lE0p0DnTF1h4qdHywgHeDEld9JBPbpoo82e5OC23TV+SuVT4hFZ
iYmMdC5LlXsTDdeDFuoN79Jmq8RefAm1+Dpe4J7uz4WYiPru1gY+4lao0CdHLvUTGSt4zHm0jrIZ
URVSgVQL9HiJmwkUfr7bY5BvWW51QyT4CYDEG7T5tSLOMBt+4NHErwjMR8uks3ZUDyg+2DlRSPAl
AOmqoFp2h29qVp53Mu+TvsTScmNGi5NCah7OoGQ5B8Js5qvQ7JyRtX896DLN/XdIUj9WS4QOrKrc
a1AfL5JRFRqAvHLHEyV6aoWY+Yu7snrGC81yS5GSj2B4HmXmO8DeNe9URMSobJC88bDXfM1sdjZ6
LZoN1zhljY7fFGYyZtFwSzp6C0XI6EupZn1wxQiC5k42dweh62DMZLCIvuOifOSkrevetl7PrySL
4Yw17IET+tNctji00g1Um45gspo5bNYC5DsLRXZJLwZGpWKo/LHPhh+lDBVFyprq0Hr1s4dzIalo
yAZdNYVlCWzpJwaD0GJobGe2yuQqi+K8dVYB6+NXiRidnb8AGopvX5tsr3Cm9MBzM21gtHIjTcd2
vk4O6d4xz3IrAZylQvg7frz9ZazFCW0mgQ6jM5yxi+muXhbhIpfK7iJZTi5pxTbbqYHDuWUQBarW
W96qYH6jyu3sj6OuBttJVMadDO4zz5rRI52lHLg5lOUZJvfeeH+wUEGvhdM0Nc3GSF3yIvE6h3pW
Vk33WISn2IjAFUr8DuNabBuiNORN6szBmyrhjeY1TyWdLTM3TzaxptY6P2yVZLS727+Nogd0NCBn
A4/F41Fr1xbP38DTgypM18iKr7gw3NLgr3h/F4BFQ4bj1nicXFuy0EwIWTpMnfhDkl1HBd9+NinF
WwMvqMl34ZQxjmbj3utgQtt3MlXDx8F1PzPgU1KRYDF7TAkmwf9rkta/Ed1vh0WMaS3WvDI/UiXe
lrJKpdWsIA3WCv1nMOTBXK7ter2RuVmOx5p6D0tgfuPAbhKquxuGVTUNKfBqXZvZd7vDP/5M2q0H
6h+3PuqZ0L897k2b5gAsfU/krrg+uD2DGFTYfpe7xq/fLbjmNa+/1BC632QNzz2LSkqqyWDHjy39
z8xZGVIakNzBRrqJq2s6xPGOkJC/p6KlFsvXagsTCeekw7F4ssqJHTeXvubhGadEn5Mc0+BXt33V
T/AuCRBqCeibJNNZkDG0I6DcuKE8mbmJdoOn31Z3NunhT2EZ/HYCZHT0+A1zrgOd+BsutXNu3t/k
uzNtoGKnvOjXoyAH7mFjXL/wf7EHuevfbot97xvxs34nTkPY3A0IKyXoQkqPeCcPJHWdS2JU0HXQ
33bzJzEz+0RviEJ1wH2/OqD0uojWqo1zXM+7PbIXfNWO6yfr4HWk4VHLtcVvUqPOjD7ImqiiSd8O
1EZJnBC3WeMqvxR9ZlmV1/DfNolDu8WsP/tX1lefYMa5nHwWf/47GTz9ZOJDgJVWPsoDKQluqWFK
YmwE/yTvcawbkL5NJg1bLhqSbPYt/SbrxZGC379c4rmKciN/cg7+Pdfo85TOp33O2vO+JrBybP2S
FrsI8nKoitjSwjGXWtBdDpXLeqAXb0N9l7JOszgI27FTWA/POJEAeuFI2xZwR8DkAA493eyq5yRu
gRPCljan1ZER9cC3A5JmqdedvVTc5O4xX6ICKNCgVDymncyGmfIg43ps9qMXvLwyGeBrk9104YR6
8PFE+nkJnSdrHarFrg/VhFiFUY/ETnbVIcmBiVC0aXkRBKLC5GolgXRz5jmPllpfBd/HEu6l+adj
pQ1qwKNj8jcXKZwvjwuHnmWKDsOoU6Rn373c0KmN3VIPmz7rDWH6Xiyg01hGgukfqp+HFR7GdK9h
LpT39KBu+a3jSLw7ETZvqBSpZCr4kfzL+G0mehPxWzhUl5uflm6m3u2LzR3X3x6yO63PrDc4V1X3
jyneNQXm6eawrsytSDaqzqQwTm+c/sJnRBCGsHjcvAN7KBCJBT66J1MCblTwhp/SFeIY3qCbDXjB
rmuL5l9MIJemOcqwzQSAVRSAnDsNdcAHWlSh2zgjIExwD2CoG0R5YHK7TGROLB45BFblHGnGOnP6
Lm0S4lZcWwqquCYxm1HOQ1C3YDT/F6W0shbBJbm72gF2qupv6sP7hPkFyEwC2E2ys65xy81pJ5Gy
Tjy29A8lngShFdbKtCKCIGwfwiBSjCexRUHz8fcViSrw5aKGn6b73h+5F9yeOtPyesJ57Q6rsgG8
Fe47GGgVIAAhCXbmMYX7J7o3faS0NZk0jNUvLoSZ9JmwVoQfhK33tmfQpTLIsGcBNOIliZZ6IR+J
2ben+e4PxpYkTZ3ualLrSRxm+rX5mJUp9t/AI+N2Rk4Gu1NB3LBCEZt6ptDMquAjzgvsAZnckWhf
mQD1wzRAiUhlnplWGkAszGXX7eDkm08IWcamCfS0j6YYKDMbSHB8NWF03MGpRof98GfQczSGGgcn
D+4zTditvEvE2VmGDzAhfmMNhM4OLhW2klEK/mvih5V8HHzMXY/IzEVNB1y1qNjuWho7RBIFHu5m
edaah9u6Oh//mvzVEnGisNc2e/9ZIWUqKQpAFq94I3M0SlLTcotcL964Kp/S32HklsXPEiUGz3rV
HGmC7TkHRVCVSoYHIL4NLMMzJquzYz+wfpWpnsx5cfE7OUbflamLbqVLGngcDpFzt9jsoy+nmBl/
wF6KdCEpwE58XECE586bFvNNFH6jE4cTRckWXxgOYWZBsl+gWN8IfO6mveEIOGCzK/7X7z7D0Sxl
C1mMSKPoGAL0t7TKlnlqeWqNV3fKuDMhk+XkNR3nHc94rYAHosocu4E4znOuqrvVr4BftFGxnm3R
K4U6qnF+HI/cTI7Mj9ODOf89bsoMDnhvYLN1wohTewC1KLP/ZuCt4XjykENZvzqSDdLBp4/qsetS
Qa2kjKGHWxWH49CJchiUOiYpTDBQFcNOspuFBPIwej/pcejzhVZ+SI69QwsrbtlNkFcQiwufV2fj
A7OKG2pxzmF0M2QWZc1rxjWLBahwHYfcvBGEUEqluJq6y0mTOYJCjVZdfDcgZNLcsZvRj+4ufzLs
X5vgmABrmTeku79ansjRC0Lda7H8fxNRKVXzhytRnPYpqf2sjTrSE+BWQSozmJmD/czZoUhVW95O
mo9U1W1H0EO+y3S/IegZJIvS8MTVUae9GC40eV21kv7QtPrAmd/soC2TYWJaFSJuD7LHIP1qVp0+
gdqnIZKMHIa5kM8vrpWR9XiqW79YtD+4837veqk4l0ajwJZsByVlpBR/5C4GGrP+z/vZDLK78IHk
JMyjeiSNvTYwFpGSA20/ZxrOQDFhPQ5Ww9XW1sa7jLrgdyxL5vVFoH6N0wVyEUG+ccFbprMRXfv6
Xg30SE358Jhrg8OgaytblsMECaFZaqAM8Qk92FnuP3AURMKYffQTEl21Dn3gq0jcjw28VA9VGqWY
gaXpXjKJ5FQsE2d4is4uRSvzaF3xwHUwaIPO/7uTlHiZYbWNtcPzuDYa1tClPNg5laigTQYV7TX+
O28a8uOZxTxdq/N/iMMeF8lDagK8oZQgH7WfTjLHk55i4miHtBDBG6qGzaUbb+qjOx6Au8f7n7qp
it5JkXpRn2z1NahcW6p/q5wVK4UoMV92T7YUg2HGXHcG0M7TJgwL6H5n1MiYSOc9xVS33a6EMbyE
GF63jTZlnpM24Vic+N4Ai69zulxfApOzLcVIM6gkdB2sqOW2sft3NLAuksEMVZN8A/lsgVVgyf4t
GCW+lhT0/R1iRTiRxQDS0KZJ42BNy32wJe3hvbS/Tl00Ph3vHXaVszpCnmx/XqQkYY/FJL7Pxi5h
Z4WT9jN0BHvL4700zWURN9Ekof4g45Hi4EJTxRyhkcGAwgKqbz++O4rbeXv1Ul/BK4ELy6GfUsnC
MRra4v99xU5FHD+tHb1p3yKWdyugr+fHWqvvNC2gDVJbNg8dwCnBTybh/4ulZRq/zaWy+Gc5+WLO
Rl7ohphEfnrnhKqH0LN4xLRpLNGAJjPx/QzMTKh3VSENi8fH476GKN8GgaATKtb7/f072VWr+isz
3OSQNCi3R/lI4N40xsy9pKnqaN6DJMn6s7LkCFbKAFS+9YGde3Uw3kVcY8iCluJa027r6lIeZr+9
BsVYDPnC5UG3zC5tg3ZnZxAYmc2FF02KjgVL3okHhOwX0Q8HTXi3EAqJmqALBRSCJmVgfxjD8liw
L0Ca4MhAvlpz9hhBNIVoPB2OWncdYfQSmmaOijGMPzy7OTd7gSVg+Twky6vHqgOMy7da0Xiqv/kH
fYCL6YkXg1hu0kbLRux1EQCxS+QNeDeKLUVzSIFP3t1obYTMudwc/NRATFe/GqibUEhKx4KehYVU
kcnng46SvkXXM4jXrE9cYjc0jvE6Gor7dki21h7t1mo/eO10loe/Hn0uSKY5z736H/t6zUfB0dlF
HhB4kC+QAFwS8OG2Vv+R3AQ6vpbFoXwvg3cyFQoExcrY9lgZITWtRUmK6WegksgvjcKxAGWjqR5T
IvwRfmBzfyQBtAminpmtAxGj/Xfz0A6ieLgXXIsbtqZ6p60QvbILXek7oKhHvyTRB6CVsD+8SoRr
1lBuxRU+Uoy/pG7lwq9oV8ryi5wOl+Lkoz0Wqs3NXBn7FaWOlgtGEpwBhXPavQMSYxnlnnWayHTK
TyYKq0Diz1hraxh/5uqH5g5GeEXIdMCFWbN8EJaj3IisljHD1JOKotlBmXcOsTQsn556997EdnBB
L8DH2XT+bWMFdcK42O0k1Fv2g4Lzy427aU8bfQfEGhEegSOMKcKelzPhE7HvNdXme4YPOlhJTvAb
JNxvWVJOjZlh9KiZoJTuh0UPW/H7ozzatyeQNxKMPpQ8qcbUuMQL6fUUqFWoP2FyW/dJ8Q7nk4da
DpRFc+FTgGXAU4hKX+uS8xDQ1c9T/i/s19N1cijKkYo2zVTX0xupGspeX1WMSssr1sSlxD6w64Na
//SKvxvUocjQShkrQfzX25gQtDysREcSOfzjhSo3ZX1tWp1erd1sUym2LVJ8FOCrkEpYO4kiDg88
yBzfQapoSe5C9aXzXb3zNh3PsdP3qy7+UzbJDS9wnRYNfXqVbcAE62WVgkIV8ArJItmm3119DftQ
MOgs0iwnoqTyliacJM7HnayyzV+HQV3gVJfqvz1pzn0ZkTXhpBaBIXtJJ/GDKzGCMiCrDPO5iFn5
MQyLnuFNYfrtq1gxTNmr26xhPF+twgQ9aZOCPBR+rXG79WhATsO1BI49enfRVhb2fVXFU51ECbNV
w05k8JnoATO4rOiMkYwtSP3+RkCe3Ysrua7rp6FTpdhM2n+XoX/qivKerEm8BDyVtl5y3yfk2/CN
Zczy7xVA7xNYWz5c4LnrOEb8fL7arU2+qfN1fqpnUFCaRAvcyYlAnOXLYNWv792/kLXpZ85j/wxF
DDYWiHTuCGtxYlCAcfNIFkrAryy+7NIFsjlKvMBkbp64EICqs0HUHGgOZj9iR/KqF8zz0p1X5W3l
GDI3hM1v9jzKTbS/L/kHmbd+wdcyFEWhqc8xa5stQpCFshSrxzvoS7oiBTBKYpJDofXkknrGb99L
dBDe0k7HRqnQ34C7L7iVQcqaoukhF61APtpdfN12orZdudeLsMfQgqoMLqAXNfP0P0Z/GQBdJXGJ
lVPiEN6c9u+2dK5YjfO0qKNqZEc6ukhHjXeUyTOAPT6p1nnM1UIzgpRXYLkXWFbYCHRLPzkaG9q1
t9IBvwXMfKxHGX3CTePQXQCk20bmX1OCXl5HWfBSk5jAmMmQlcWv1ZVtFJysGJnIMU+ZeNCdNnIs
wMi3EdxjcC0XS+n9jP04B0JFIfexpuiYK03duwTnbHZkCQx+sFQ4zmhxxK6pe1IdTw5gOtyeUx9r
b14CENz2CiDsxbOWYaN7ES5P/GEWk3+xlTQUkqRClPm3zXjbhQHAIzudC2StIxu7JHwWUnTSZj1Y
HIiauFRfQcMlXry3yHhpfClDxpki2CutzUn2NPEFxdZPafNw8heipfZiIjzgFfK6TwT+ysmmcmbG
ZDtDdXTRqdJQWJjAXzwLullcVcCmBMx1f3exyj/jCVffs/9/PWy9kzt9Amnf06UnfVFIBIbYxoCW
ttqUKXSIQeZk0qdk9EdLl1kkbLDWeJJhxlzb+ZrlLtA1UHtyWQDlSQJUh7XEfcDRHfBGX8oI5JnU
zzdQH8d72t4DkPhfjOD1qayNnoUfqvTNJLpi3qR7PjxovZIJpNl91ax3pYVQhWdu1fZEAB4abFtN
yT2uLi609s3sjQ4ACYBJRlSTZVOmSk1RdZY7lw8n+hZvttVVLkH8Zrqt5ZEcklVoheWJuJ32ZW2y
bJlqGGq2W6pox8uEYuDPRuuia79jeBW+KDmweEJycMKmPZnkBeaiVjiilKqFfGNW5eJ+zaXpvVfv
v4SxFYJNH0fT9jbGr34ACcdhzvObj2OM9hkreWCtTO/V5vCbGDCx4xk+QMNEz9/G7RX6RtCQgJGH
Xmkk8vJpo752PM74UpVEzoGJd4yn9rAp729iRsHGCNmJiLxVcXBQm4c4qai6sLrikxj0C+cuR7vO
O28wV3rS0wWJW6SVqWYGOloGRdSmubGVDFI9cfwbLycrFhrGec5OrVXVD3zUd3bsN4iUmNRT0hyq
hU1ZJr+NwiKOcwg1p1VuVfn5bPZYShUFC3LVh46WmbMptMKCMYvdsNQJHYiqbbx9wFG5QVqHILah
RZMCLohacqO654/4Xq0JCrkR90lLO7Qx58tcyl5+bMCZQFLF2ih75FXgsVuBgVmFITrHvfYXCp6r
KKYfTiBaZgH1WI38YMHCXDLUhTnXG9tEw5ht8SgN9dfGrwuLk2urVr2XNR7xNILFpnwmq4speQNa
9N/pPPG+W9WB4j4zZUTdtm1bGRnHkXtsKb7WDN/aKjGgrCQlm84ssnXLd0UwmW7NL8Vp0OYbenIK
hoAAtVNacJq/2qDIs5CR1tbm3HldawXtViVL/ck7WmRmxGzw3Tpi3HMnZFoALdIovvq+9xaWyJNP
ei3FN+ktREKANI44SBF1fpi08ty/d0aDbMVA2It3vcZkBB0P7Nxh2v84mg0gXsqbrO3RvaESZvPf
MYXuyn/ToiqXDpOaF4qssw0TNZ+WVcSmkrRKaaMW/oBOuMbetOb92MDbxjvw549/3OfbqX3Dt3iL
Ex/EXTnqXrYkweVAbb16tRQDpLHLCru1adAX1pryUyLyW8pybPvW4bDfHKO7k7p898YzjggcbCqZ
6WFweRfzb5x35nt++uStUizuF0AfWFie1BwMELsRS/4R1/UKJhjo2wYrEKai7Pln9h5M9GyG3h9o
JzViwL12MyRB/ZWSlgljAM5z714gwM7KO2ATuYPUsndDG7je3Cp8POVxbNGJly9XYz4xNK3dW+5P
KW0ONFYWlq+8wmmsxJo04i9kUOB2Wp49dwO9/uQ0XT/sINXxpJzDMik4O6GFO0HGB0KO87Xk+n5D
Z5fcHZUlVU/suplm9Xp7od2+JdC1IuTnNtbJjIZGYOMuBG7u1fkYfcsGT4eyLsxhwCpIBBkY3bPA
s2aZCyC5sdK/HeaKhgUk0uwwPWyIkA4ljQAsAIC17JJ/bKNT3Dmv60OvOqFBrugtdYn5J1gyPpQl
AkJtT/e8Q9NOzg5l+cbV/ut3rCYEA7WgeEimOCAoy6JXGgGR2Ge4v92TdV4ezaSUWcDXR8U0Kmgv
Vd85NVmymvmD7LLnScTTAUvURdEm9PWQHIVwfOYcy3oNZ4EvEOpkTBRaXj4N0uJNnyrMGcHAcPTP
GA2pT4sywICxqkAJChIYzH6x51rwaPAuuyuUj7TdH8Rk7LRvNPNM+JYlAxDvsDPHW25Fj2uDD7Dh
IiH0qUKoxmpkSW4TlZvVmDxeIFd+s4jEIDmWTjMaGBbk0uqF8RoUgbu8oVtw0qyUwLp7LjdwtoEX
l+K71b8FX28Whys2mdpggaz7YGQ5K1Alx/7JDAvx+RX/zBmF2EkC3LvgMZm5/z+4hco9q+KPGWl+
yrUty3Hjr/yByhGCfK4KS+kFJH2xT9PXL5jw8UineYtlmtJvWx3EHe3S7oM0oQE8e+sDiobkNiz7
VzqnIH3WVBChsWl2IyePmFoz7gDUsORr5UGRJ+ri5UqD8jaDYonG52J5tDtXKLTFec+Pw5DOwkQ4
NjRJQFpDuHSx8sdxQt2m81S71iO1Zlznd+KFaKqIWgyal3PlIQu8EV14kuUexnPdqMioUMJBfGUf
IKOLpV38fmLgF+RlFWlJDgdCR+oP4n++IN2C7KAP2T51FVgerTyrVmrGfg5R9ZZdXoDcYd0/FqpM
KL6bPrZ83pYovcOIQaw96oE87smE9QRtFY/UQvzSaaRUuXe7fRe+Wv+hiRoFgBVAsyB6XC/YIwq5
/AyWSp2z8uWuY+R2I9wIYOgK43Sm3pwGApVBfZ12PTykZ6z03op0eROBMQ8nmMUu1gWigA8H6G5M
I5TslMqsjRJPGr2VvlZHsCUNFWT8UiF/D2OlHJke9T4nMvROO8cu5UHwCcdxffv/EsDBJUDWjqUx
YgGVCuXuogGEJ4LxuCbqgR0iQCssfL0QHOtBAz3OmoTTUPflMSbZNbt995WJgtawMNUS2ONJjeBE
3Bd/wdoG6ke05NJiZODBuWdu3PMhl1yFX8OuAJkSSExMaj8eHDIWF8rS1h299rzObPIlofa2Ct9A
FnraoHyuGM9az8qskUEYPAnAg+TG3sy56uOKJFDDm7jl0pXTGHin4v2CedYrY2tFF9+K/ANTyjf+
3y+e9YF9Htoq336HVf04tLtjqB6XuXmVSiO61mnaHnTtfMyOiUKAYgYYFubHCWC93/HmxgaOIpzW
OIUdi4Crcnk0jk+G6R3AMAapAfuLJH1gYNt/FLijT3aOwycgwWtuh1DjQi0iN0buaYVYp7T3ZM8X
lW/vBNtAJ+YF5qShxNs4b7s+G5fdbkpHttEfuuq2rZt1alX5y4OGDeHUfR+ATHvmf+f5eIiUD0IK
4QhNubclOsVpq8fbGfkBsuqwPpktpgS6TA4fkdfTO+Dsosu7+UwiuaEbkhWhraymkJ0R02QBi15k
+mW8d48sMyeBEUgYPt3B9Gx61GadtwiSz1/IiFq78VaLMnO5dCCuZtoNtDs+ngZ6DA1yTGEIWyH6
HI8FOGUhNAV5bPSt1q0Sh8vE4ENHxisiQ7iD62uf/NtUai2lHLf7NmhVgjrFBsib8Day918Cs3pt
01KN8i8eyGNmH+Vwp47aSBe5+RuWsY0xoP5tzkKpNeGD5QWBuz8X1Eey2Av4ZhVpbZ0TWGrLBWAl
gPb/boPl4sBUQ/p7VFJmz3RnlPK6hfOfwW4q+i9DS24dnv41EUeRpEx4LVT5OYUZOQRzDtQ86s64
ZiGaNBEPxWpiFpT9eH1Wouv3LgiGGmiX0VbnQX0Dv6CGchopUYWSnm8Inj6V1ih5rDhbjhEVi4vA
71lq8qfIhJRI/snx60LuDQBOzMjWn8GJdfIFZJoHJU+r+lbgzYsbiGW4rJP15RQAnvFOZYyhxtXg
f74yxU2/L7bLKvvJInguQJ8b8W15KAJLNOYTebBWMH/cYbhYbo2nBldDO2QH6IekwsejEQPO02Dj
y35LTkyzLl06NfVMzANOEhNKG++bAJZ83ysuyAUdrzj+kGscWEUjXcQ4Vz91yZ6kXBLSBepXHrAS
NwOpM30O+dC6AB9HZMMssD5FgUqPcOyRk5JChQmh6B5Ble3P9jEj+7WVQNCgDAjpIncuL8iUvHM1
FYV7UzO8+LZbmC+qoPW1kGgKF8aB+o8RUGk45X9e71Li3VhH6wDSCiJ82HqWpeAr8dDKjvE44w4z
HlFh/bHnctcpQ0fZAAQuLfx8o9GJG95W9yVZBTUNgqEwQzBteOFfl4ZCNaB9+zqNK1hpgu03WJ6O
K1gKDxNUax4JJBR/jiUcuK2ja8jCLXDBonVw7XCR5j6V6w8TOU1UYrSZ/+5Iox6e2w4syiX68FKO
GwuAmUYfwX4+J0lRp6q2tVIRnnAcWyQiWkR8EJFTjWWLlGahNuzGkV8xKC8yq9q69uDtjVpE8kED
+H4wdvBiNL5UWfk9APKprE7/ZcErBCKe5coQf0Pvea8Iuqib5FnAClpKjqoJToAFVEcGTzh1T2uJ
240zxlAR2yj/gT/tteepfVQKaylpu0UKe0szgxEDM9HlWWt3hahNb+j5so6TYbK966cXnnB7lH3q
qSn4GLi23XHghBqqdDn9toVVN8mzXmN09kYeOv3Y301nO8qNnw46EJmO+IHnvDqUt6M9FH/T2Fzb
wMy2JRTVTfQT0Igika55CBzjeMzyVDddnrRZNaXC9z+VHh4fijsE9m9XL5DpaFBZwIeNNK7wOrj9
5XefrrTbauiYCAZ/QQiy/7kQarQShs6/DntfdvTiJMLmAIqAFV+4Hdbkgi9aFOmeLyGZheVGcMwg
EnGy6eTHjTDxiTgXpZzR5oSJY9sge1vjvlPeb30TSdbRfw6z/IUcH18GNQsyLNvcIteyvhBreIJr
Naoyk+ao4sqEMOFY/eKaaEEOrsx+bz9Aekb4I1KX0hkGYa847u+4V9pzwtcprXS/GIhRoJzthjTo
2JVzSC4BbZJfh9S8Sh4aegcc7UTTkFWyY9Yagmcs16bdjkVpyopSoO4aGBnuvPMfO58JV1ZM3X0L
dvALt88AuZQQ+TSmlPgGWtLMjF85k/4xWfTeq1O1h8UOmPxzh2dep4YcoxY2m4RyfezDLrD7+9UO
QEsa43ZzurOQt50TWK4m0mIvNdpXh6I9bm4IpI/iWkAD4Noc2CnSLppuUuyKN9pmWQpSGPSuwUnY
2MtzsAfmXjgPBA6H35gCxU8nH4quRSxxdtvRBlSYDDs0lv55XByemC+T3t2iu2pwzEX1BhHx/mln
2QSCww4LV6GiKpGPAcdCmKOuNTGFphQa+KdZmrQJvp/ftHt1noROOigQrnAD0Ow/0h/93sI0VXAm
d58i2LSbWPDyEtdfBlHswbY3Ysa3HHBVsBpMsaIg10p4BvJBs103W2FyCPaQswpqXhLmah6yuVq6
ccF0t3ifypG88Vpj/Lpcn4WOwpKMOMIG9FC+v1VhpcRzWcWoU7k4u2gHVoKtYPUoGnlrMGuek9/4
287CbLIZA70j8phgEm+X5rIGLzFlxw82aKgKPJGdFUPMotyChDURVI7sj1Nea1U0NzXvoCDepCX9
jGhDDJr4pq8T6VyqDN8H5wePZ3tHdEDt/yxWp8dEcuBUXmwjKF2r7KFKnIvisb935vKwUs/KLxwD
jPJNPRP/vlVULp9YSofBu4XO3BcgT/mJeOIHftOUw4CmC9HqxNH3q9uzYxYs4W6icYhti03YUqDf
O74QIvjiryuDZyMCUCUOV4kuDHznb/b8dNgGEtDmIuKmRKY5qmvrscu8WCDf+u8hReW1ju9LLNqb
9GNJ/XnzqalEHhwn0JS9vgNf3E0Dljty1GTyKNc2feFY5XMIBZQb1vxAcX9gfPY6Pa7CNKpHZ4AT
0O2PSxe0onNbn6KdWYpJr4uZ9UDoTQSuiin1OwYOL4TUOp2YDlWIy4byaYiMqcoIoiEtO4DMpvVu
x20TRmlJ09HTORK8Hzyo30jQBPpW1BQBmQzQCyaNnZtK4+O0fXMsNDohKMJ8yYc1xnLaCX6cHj3f
t0EwACdCNncnoCicdO6tpGN4f6ovsu1smlz6CLc3scSEGITwhu/kYPUUjrF9JSl4/GonWdimxfcx
88aDZ4bmfiH5EuEz7Re2MqxAkyccDdt/zeOQ9NeR25FoQCnOmav/t5d52Xs4VaHFBcaruUctncdN
+IhUwWLrIGRZz/qQ+xKlrqifJxWbxOTVJa3TY7yK1ljaKfckH5Du1Mk6fMrUf6EsDdUGIYz1SmXU
K+olRAAAFwfhsasF37MjeBjbbsSatIajc+DJ4M9Bsj2fATd/CJcqI7RXbrswE7ZkeibIGRXTFsDS
M2h6kHhRNHbIKiDD/74gDKe08DgzOv1tMEiUmG9P3zzgIMU8EMZhCa3eiY/tj/B+UQbhDhZ6axni
zm27GmSFkwZ3TwGz7h4/jCIhU8NQX7ah5XKR3Bh5AKevTLCkflr51FqIEt+FSxVTM2SWRbvUuMzA
Ty3aPG9hlUlFXBAWQO/oFVsO5wl+1PkCPzIU/KnJnBiKyX/8hp/k8wSsoSHmy3YHgHHixCSYTfTE
emZWAzodUfgglB+Ybzx+YSYubevywgUcDpvMrLyLoZqvScntBb+kAeteM/i1apcjb3C3TmFoVhA8
sSgulAWmmjuE60RFYoUGPY8rPJiSc7Wa9Pta+g6Ck0Z16ebHQPObz4SF7vEeggHUplFpf7QCGAxD
QCctCABWpzsPf0LxYL1ydcN4WuZ+T8o1dfpZR6yC4LXyg499qFuSGVTHUyWH8qvoOJUrxob9zomm
fP7VbXIv4qzGKVrQDTIW5xwABfHwfHaudgA5Udivt+/dT79mdhw+JLXVnpShkV4YkwO2NfWV4R8c
M+ua9uUVIRj/jmKbpLOFk7iYmepjfvi9pTQC04diqCoqopvloJIthkuL+AjJ+nEs4SUcfEoBmlcu
TR9GKsWD2QMntJmLFVgX+RmjWxEW/Vsn0KuMaLhfr0phImfdEkoZBKHHuTarewFhMuFqzjvE9xhm
cJA6khxUegJMXC6A3yeru7RndNimMxymnVR3q+JF5a2VjFE5e5yk5ozvb1c8io10xYTWVyzkC3bG
+lQDSCu6iA8qOG+0RR9d2z1shT8WCJ0TPn0+7m0CidBXVTvHe0gCfUIccGjDoB7JjozCxQ2Vz7CD
X2qAAD2STUehsxtK7atMzB4SCit+QufKfiZrZ5lHWXO787q4CRWUX+uuRiQQSmxNOtoKoMVUjuvH
VUQYGU28ke7r8RqCQczoILSvQE4SGnqhgYJgcoiz85O89PJwVOF9AyJ9BLE7Ff/vq7Vi+GZpNQwO
GMqmEVV40j4rmkN1g673tMZZTIZzFTwdVwQMtncLS/Nj9ep5CvnZeo8rmnrq3aGoHF1FZKqZeA49
fJbpQOZfaf4mnRYKnvShGrWOrwQHdeg5b6wB0IQK0R4C93KyuGLpzqHc8Xl6EMVVtxJqpCAqeSsv
64AcJIGYDgLlQm35PoYK/gD+8wxIWyRFTAkJbxVv5k2kM0QlvxHN/7zmamsm8QM7S1C0p3qI2GrY
zVL2BHMPOwnOLZB6pifpIDb/oStlNjcdFB7UmYzj1D3RDdC7aiDK1NvIDtR4smnFdVDa3D5Q5/qB
U2kW9xNZbVBqz7l44CPhvEXeyXbEJx8hQuq9rUv8C6yUQT6ma76tNEIgdRHC1z4mZlit6c07Dj5D
1HAbSdGbiVBpWe9O6nLO7ao0GzWVmMCM5pf4AHTnAlHFevvuQqXXNlKo+586sawfoeLNZYXys2S1
nsnib7dBcbS73Y43jOk8lzbDa2lYO4UnuQ1S5Z1w5fzlngdvBOkI9Lj3kywzkAeEu0bZ7agF8eIu
YcRwS6JVeBL6HFWCco2hsPf4Lq6f7FIN0sYGW0sC4wBRjdM2zxDXs0lLKtoszvxzX5JUbJh6kLlT
nvHbfB3b1hzU6ukkMvKH1V4DNELPmuLiG/GoGR3Nw0601eUBxtVH5084Rd+QVLUh5XIo7/PDUrK+
+5qXt6IQm6SlW77sslwMQi4xPbexDvf6hGbjHo9tyL256TzZEtstZu7G3AraLtgMIodXLNTYOFlU
Ogo/2eoPXZCWVYVrw14l2e11laQVkEpEboNuA9ntIsZQxQENv5duRazrgLfkWEzeK6MzQ/CqiWqJ
pMDMz5GdHVDHsOQu3t4bf8Ztn1Wf0yShd5or/ORm5/y8pHrtMk18O6J6/ZTxJfOMO1mOXJMTRwxR
86y1Q41qbEQ4EbLJzAJQEtT8PybeV6rofzgvBxIg/FRGU9zSN0P3E/zmTLNnOut7iBNYKY0X0BU8
I1OBnihNQdICHQYjc/i0ggv1KnscRBLRAz7JLTPPl3lF5sND8fxY75vmjPBeOsyeVx46OJ2osK12
NUPENgq/v08avSbi6CqO++hWb5ofn6k2X23QfdsUVshV8vj3E5O6NhSGNXuKV7pNvqiuUzaZ9Dq5
iQEbNKq9KjIgKrGR0tvIdnpMS7DoJVq++eUV/S/e9TO6fMqE/TZ6qBZZ9lf9s/oRGSDXWd1os5Rx
/hDiAjOY4SaoXkv/lcPwdbmENE7WTMoDXu2q8v2srxWCkNfMt42dJ1QOMRXFMmxgiV/KFdHFMBeX
JvDsB563Qzmqu7itf2uJi+YYWDL1TLczZsXpk6YWumlPWiOo6KcdMg49n4gvF0NlOVcvZ3nA55Si
TaB+e8TUKYT5Ra7m08Akc+zx88qhvcD4+8kaameuek6yXLwergC4PYsNSBiregCM48QJzu0w11pk
1S7wt3yo1bTe8J6NLnxOTGbSiR7EJ1N87f1RQ0kUMeJanBBEklm8UpwuMC1uCtRkdJ5KKnni8GUd
ehj3q0I4YA9NmgRqrHsIow1NfKPi4vjzEyaUQLnD4TItaF8vNNUFUR8jEymG+E/GkMSnXVgLW4oy
jUuagNfvnztrjZumy3Wgtsjr5+PLefafpC9aYdenrsdBVuogPOP137ZvEkOy0KbVypp6Rb4u1Xe1
ojzr22z1qNggEHa8NcYl3ay3CRTbGNKI9LR6z1iN+V6u0b+dqU1mZmrjGXBKUAjWjppYSIGWlALO
zmoAocaUu4JL7vwF7yGGHC2RUzx1kNhfS1VmTSamJ3HDc92Pc6YF9mlskF9z2GA3Yc4UNREOAao5
wintdXwiSszB1Aw62h3bXinYAUxEfme2XdrRe8RI+MlZ8fvuNprGoZJCg3AnizNiR+nS01KlImHe
jOKejD5+gawUpXetcUE1uerGXg2nRr2+ntO/TsL7jMIvPTbMQ8YoUu4ad6+x9hXM2P3+CK6Uc1aV
Cw3BYON4OqYgUYPwl2i+KnDREuuH/V4ZWhS0BwtYFQEdSZDXe3ixosDfYIBfCzN1d8TmAlaDOpgj
xHn16f32kG8eALagNWHVVCPjlaslWWzPIv67V4Fr963FfCYwXs/hlvG3n8vvED1aVXGa99e6Arfo
e8dWsfA106xC0MPY94Z9DY/TPrbrKE0x4bSNaBRBgN3R2chWInUhis0fcIiNBudZZ/rFz5HhCgsF
WSOB2f6LYLq6gMTE0alW4whvZkLbeolMh5gYymHzKLezqEERZRIARnu+otlLZk5bAmiEaK/dryWq
AEiRqNU6JzVaLCFidl//gW/EDdUv7Ztun8pD7+lovuJDjoof/DCvLC2+teU7Eka0LCdSfSGfhc2y
Dd4zQm4OVXRbthKLJLKEPhAU6kavCCC0stYDfRa/p7ZSTEIYhGI1SFyqvr7ksfZqJVpiAiQT5ghw
1muBFc6UJmQeDZkv7rJ2aLHgquKGkJzrgVRC21ybAhnecP0oAqQFPpvpxUQwvp1vXL//nETzdELm
GK/3mpx1P2aXKIOTMh6pv6fkvultUv0np55yehRFsjH0cUeG39vBO9s2zbkWFW2FPgWUYZl0upKp
LCqtC4gLZMcHMIVGUok0hbFBYplJn5+K6rFA8VQmixenkUYXxiDnltj7f/7/Xd9eTMg3DXg4ribJ
bFk0Et3QSniHVOB5jkNlhnnkuf6kNAbKVgyI4XWEgjzbJ+2nlBdM/RwLLTaMX08/nhPMchuHFNDt
3bJt5UVNyyQsN41w+9rSTpg2NKMkqZ8zJatezFMCvN24ePU8wrvqt6ENq8z4LGJqQqnmrIIgN7pY
H3qt6PyO04dut8yyWgDDMBc/Z0n9h4+LBxN+EuelqCdh7Pc0AekDtNrpSH1ZIjXxHY7YNe4gAt1h
eiNcpiGgOP355Xi3mOogiXHRQW9koCvGT3e6BHIprg5j/tMtLdqzNhiU8uuehpesJhgDQOTeiYbx
FXLZ/0o/DAgQDFZU5FT5r9vbHWr+3BijCqSQkgA9lwfsAORfye4URdvf0O4Vlax0AyrFIYYnX3hv
OgaIeP/wcx8U6rLw1pxGr84uoCNtbvUCjddzNu6wJRS5TInHIn273kI9dSBzlo6BRF6tWJ9XCOeR
yPguku9zxHsgGjHRWEeoY3Qlqlfg7MgXxruw6nMA+yLJRjRLILt+EpUXlyh5eKQNGl3SBkoGOwZT
Lvi0Of80pqFIq703iEEwff8xfcmTy+TVvIN/dQQ3ZTItf5hciwt3FoHvwPJ7C9aJzkNnMqlC26+t
9INUgLzQbISICWddCbp3KRzCMNYzhgH6fsr2uHr5Fu3terXdb2vtfsy2sTeRHSjOsaCEz9yYbbFU
C7fl7zSUpmN/OyDr0wTiE4kppe8ectgHw/aZ2E7aLIqP5iHBFJ5BcdJMbdD1PI15rZ8+5AEv6qPq
zMk4Dt8jTF7eYh1XqQI2CIB4dGWshOqIAGL663y25U64+RNM3YjQUzuNSdl3Kr3U7m4cKQLlLCQD
oh+1YVNxE7uioT3te2US0m8yya4qmO6Kgucv3tpYpqRXj31imwucbLbvYtiILyLPqIBwn/qMVDZ6
S8aNI+H4TsLFYLzEPp+J46PVYPKkMb1lDKwrIosPpBMSJlKtBOQgLAZSJYyuxswNZ4/DqUrR9lqw
mEyF0xp9gb4Domxde/LtQKhldwQRnslc1KzleVWq9bbZc4GoNBwLq194Z95Iq1SuL6IeHxGu6dwS
xapBeTSXDEwp5MlP3rj3ZZdVjW+pnImLD/gngT+/3QYgOmRO9p5dx1hO9tPBarNR3k1FPuUxiOG1
EUc72B0ruIsQM+nY5V15t91g8l9ou8O82cToN7a5JAlqgpLGZaJkMxs0iAMSLik5SQMmf8Qrzc8g
MUKUu8drWiYL516HboiHk2vQY1ue/Hf9HlmeIjPvjvjv/q2aPXXfAeHL3+w5tsBowuSOt76vmXkG
HiSyQxOCNkmsRm59KPYJiwZSJVpuLnmSr3sNB3RHvlhmmSE4zZ64vbOfQ0WNVfuO/cSvddHDH1uu
lQesxtQ9dkglf+TpLz7UJl/2sTTugk8jscBvAZH3Q08nfwlob/O6vHhLHcUcsrj0Xz9zsw1T7C3R
TPINfv3Pjbivw4EISVo+B/WYKbb4W8eYub3lto65r0UkDB8wFyFW33sQeObLL/M5sUV7/6M8Q6Qq
Hr4RzgwTnTaPhRnmm+XgMx8gc9f4gAIvTsGUWoVktH9enojqAiPtYHclxyzlhqB7Zmwx+UqNBhfO
IoD4UcTdP0FdF/krKEA7tl5WoHLRjwlngtWSKucRCS7y9qSzJ68nktq+c7EGNnCfGbYEyrfIzrUg
mUOdWD92EG1wtPTAKEPS+B1BFISVK7GiOWxuuhlSQX5dxU5PV1qW+cxbJl1QcQ3e78JjXTBpLuS1
BiaYVsY2QLXuq/zTK3aL3gl/4tD8XeYT46sG0Q21PIf8jpXqLvHqYk2TDjdv7fMZkVrtCvmf1P9d
DP7u4qa6SrMSYQqfKPcpqcY4TleC9KKSXnme+2DjsHNKFeiU9ppI+H2IcPpM0b5PTzGWotxZaoSS
Qa3AToe+Xx6rH8bkQz/LdO0l5TO61Joou3WnwSrPdXWIDKYMAcWpPfn68iksToZUo4H5UbxUnc2E
jdbcQcF1iEG9NIrW8ibPKyUfwciag2LFzoKf/cd3RBt7yOCyBuW2EHTMxBOKIhlNbw+4fNN91a3H
A/w/7FRMmZqpp0GEMIva3nBQeg+7W91UMQUjGDuaTQM7UAdM6F/FVt1oZwxmO9nJfO9sUqS1ocAc
ERQXoM9BZx+I8auL55LD/aasgWDca1n2ipwdBooFM+xZCM6PkErATOq1TzO5EgDEoMYiCk2U08vs
0optL+6Qo6ToXZOgpwBwbrt6L/w2mfl7LXUlS4tJ6+dy8sL+3Rh2XNtPWk5Wtlvlkt3wrVcVdWCT
npbdE6MNCd7ESuuNF++gKGfmd8MwNPSiEjZLLNvai0dYk1WVpyWsBikU1iKizupJBIJV4FrSM3kT
Y3MdoOKVtfRWyziMLwgug1XwbTk1c5Sj1yeeKYN5n7rP1fTbYq2gJEIoHOmbVVvca9HIJG+dPwkM
+2DYxJ2yzItKpdiB53ok0Tfq3gaokGaeSOqNg0xDU5lX4dandZabyz+QulWWQY+/oy9CV5vpVbe8
s+9jE/L3lOTN0Zrskcmtlwz4FM8NNTq4S/pRnxWeSBCBNJf5KyDwVrn9UZUUbX1T8YyHZqqBx9K5
TZtpCwTxUxOp0Pr8yG4L4gvnSXFS8l4ERM/9FV8TMM0kBbenCU/hf79Li8Yv4JfDR1wxxVfqeV+v
5uaWIteWgeudtYhrk0emuVVohJSqHpqu/TmpmXHWuOt5SJ4IJ48BmLir7bQpwSjH5QNh+ET5ZS2u
+4iC15K3PWlFSRNJSNUSTkz+YmEFVrMPGFhs6zA+i58ZyPdsnD34EAbZEmCFTzAdRAcOg0/E8OTp
B9cSWJjcNWecOCZD617poT3dFnqsHz9xdVsoI33V0/PXMWT7FnmEanpDUf5Q9v+4SOwkJOIUj/U7
lSL6UddIJjWdeLMrs9NuPgqU0xDodq9lN6Gjua8BEutqRV6gQK+i+QE+XsRFk8s+g8BPYwnqEXC4
CE5Wxs1AVpQdKSAEnziCJqriw46GRVPlFmvUO+seSk1yg8fYYVyYQlzuqGNUdAi/wIroCFkrurhC
KM6zFR8hqZTggCiFaq70r3dRsqdrDuj5pH7bi5gF/WSwoB2Qln0J/71AQ8l5KMfF918weKcaPCYJ
HCi7TDT46s7Q3tl8mg7g7I+m9ur069M8ezjQeKFNYYwV13L1pkSMXtRYH1Zk4peU8i971Ft+RWzh
TlMw6KaqEhQ9awm+wmHMdB052OYoUiXwSyGj+EOOXVGVOyCbmUgqSe7PHjl8nIiLGCivI57OmHVw
2Mlue8IQLHeMEKh6j3WbeIPy+Dib8FdU5QKnHpjMwsmoPbkWinzJ11nbmgYBA3pedCsCRRwpf6ZB
6oNYT4dLSTOHt4/Yx/jUjuHfEpzxmc0WJ9iXqaVP7v+4zHbY6zMm9CZmmaKnp3ZPuLiZQayBKTqv
4NnfSr7+B9bqMltnuDn7mTydb8tTlg5kKYQAiEQcTj94lePPKear9fBNi3svl7E5j9e7f3i2LVhz
rnJxy62f2nfwAkD5GAZb3o9jkOQO4bXt2EhE/K14IXL2Al+ccGkMr9NIZZhfPUD781iB9TfDemSk
LHz6F9DqN+crPWOdMHxwOUKrJc/Z+guZz8FIsSjtkHZoMw+7ycRdBXOu5+ze2c36tB6Mq0RMW+vV
wxEPnVtx9atM9/ZLPsLofQTem5AHMujTNhiXitgJTfSN8w1KBVTAthhwoR0rPtK7N9PxHW4LbuKG
AobCjTKR8Uv22RkSLLsH758YMS2PXnQVhR9zRC1dVrmagAKei2D0DzAax2E3jyWuxsMWBD1nT34n
bxgOzjtmu2dU9SjYEgozTVKhD/VMjZ3UJQ9CbJ8Qt9CH/9cUpeAwPwgp/6YNRNOfdHQbxVAuZ3XN
GbAiZ2WRo0ytoFsu3SNQklHP4e4urVOsdsh4tL9H2VQPNoDLPT/6JebvLPrPPmtp/uTciY2dOJmN
+M1/P5SWEfyO8xR3SjAWSsPjVP+URyPOkOg4zW2lWfkXNOdRICqPtqhmF9PM897JdUlyTgzXf88L
01T7ryv5D+Kyf1E+BsNHjGENN2+VG5yPBX90FzqlojBvdccCNXpEQ8eidEhtyyLFiH1WFfqc1CF8
Rk5tQrq2PI8YvPJ/SfReoJdyKQ8yPK8nVBZihEt8x/33lE5dwSBL1HkTMWZJ4DKR5rv8OXCnpSfz
w1q+unIcowYQarjZ0GysAc+pzXp6tUDf0p4sR/hzwTGj6gCIV/cmdRmu2zrbodWJDCr5sQ57tD2X
460ILkGSKZ5nxTNi1bYHwP7QVMywJNiBD5EqE0ZFDYADqxCsNBzYUYFRHJpfBKuGpeUzsUmYXv9L
OpRCyJ7dmAt2yjyETS+cQ1dZZ6If0HUoS/q51SOjy8/jbhCpEWPtQbJF+u4We7MN7QhUf6bBHb91
eIbqXkbp56PvHjCC3VMG8eTYEgk8lF8VR+qebdMHHF1WjJq6cWGNm4RsjopU45uIyPNNROxp3KFt
9PWBMBj6j67p/TRWJPuzMNuuXAvH7WdOArYPaD+AgHhGkFNFJAboFSvZH51h1DkDr23kkTQIqPPd
E530jiEgHCSeSAt8j3by6qqevGTWolXisa0mL2VqDq/knIF7fE65iX3JnDy/PU826KdCSseLKa0U
0pvDZTnFjD1zOZGfiI++EEF39d3+lnDhD5zaJF4VC+tZ4ooYZ9lABSv95bV+ubEAGwLZQKHbnWLX
7h3YLWqoalLoFfV3v1d6Y96ZIhn5GpxtIEfxN+ZiN5ZT2yuR+WS9+xmEx+qMG1vWRQWGUAH4w2AG
2Dd7drj4kxGwyPgnL8iP9eZ0RArd7gzqJyfAL+pGWjgKgcp4UolXaNuYbYTCkA/5uCUoouAKgtb+
yh4Ca+3a1tm1cBk+kMQAafR6XcH8QgdMtxA+0VzXkmcQeZPntR1KLDErFJNjNmkTmiPsDuKZNWWY
4AgDSXB8M6fByb1YhnyQaaOXBfQeassSgbdShHy4/aAtyREl9p4CtPu/EAb5iOWVBakoM3RJj5V1
ZNCSsc/MF0FEPvnZ9cYNt6zcIUz8/T2m+wcZ03WZ+5tOrqzMadpZMn1ViO5q7bLHDHpTOQtUzxeX
xiuD66zyP4SWrvWwjgQGAKrvsHwgsPecWd3hMKiDHsU1tAikqZv37YufcHMu+UQez5Y8vXmN9WRy
kJLqkm4bCra752iuyBiKlk8zcB/1lqudWOhf/GDvggeG9zCzA6+sYazldSZk1gRHsIRdmOuEieTd
/ZW2Ax93lyLyTc/7rDaxYirQ3HDBpVzIOVkdd8t9z9Ytiu5dhJu7DIPwvdB/5+ZNG4NlFzCYCkwq
Fe1GNOvCzGaWXMKQbhoBzxU8UFOptcErWLOmVwWhoN0+CY9VXABtF47zg6pNTr5PGgQiWPnumQBx
cHRKjzXsp3eRhv/+xLUZ0y447dJtNkBDyxqGdR7LITFexpPlOxOyuvm8ElE360RYtLaOP1wbzF0f
jps4j04blkqJpW9vj0lxFz65sdiA0y3yjECsswgiVHSjb1lYnf+gTDpEQNLkVWBAP55cXqH/mzWj
uohIO++fyRmAkviCWtLddHPpDWa9IUk3MBOlW+9cykw3vjVf95c9jx6bc/P0KebVSSZaCsGceubl
Z1TzBAbTwX0OwNd8tjYudDw0otp2rqAnfxPhsp2dTvTt88BkUc9RAV8ZJJtwgQtm435sXHqmu59C
7wYE3mPqXGp9QuoLHt1tjPRCNQekN9/575HdNsnmXQ5QSDS2OZzcCdmCBPt/VOg9umNtHbPzN83L
M2BAAyw+f3rNbibOuOxdqS/85pyBElatWo4vPi+PuBiPhoRcbwZ8L+tIvFmabqQKwNqv8hHO3TJ1
ZNBaqt+RetoTsMleqEuHE1twpSW1zHbzLxL4odjyf4E8zhRJBZm6noXN5bhI+HKSgpOKKPXhIbk7
I5OmQYPf+YlasHhHpWnTGXI7kzhzduvNkEDTBHxrY056thZABek6D+id1lryVJBVo8n62s0jb0T1
sIk+AwL4Q3CdoV2BNHrXO1ijb2LnyzJ58G4C9dvQYURLhcVwYLUnZBF+vQB1T0RuO6RsqS3hUs3k
QYWfrg0s0j4TrvVPszuDz9Sv91usO2VzeL5Pt8xxiTZbE5xI8tLBLRz+FW7l+mJGQwf3nPu73Vmn
U7vYNH8tDU7zNyKSgrgAo5BCcnKDLjkzL4EITw/yOWAEogd7vxDtfsVUSQ5A0dxnxKVD0z63wLKO
3GP9W8NtCdYoHlFpq7ZbSxw2ZmzmhouU/xI12QSIs5WxcqIb6FSylkJLXgaP8oEpmvQ/hX50x64R
t8nEGuQYHnT3G9YUPcszyx4pYrsephp1QHEKGerakjlCeoY0yUx1rtbnGZhC+tL5z0H8x36CvOJX
Re3DGF3DQT7LahiWkW2cJbdcJI2KFXoADxvmNK1XKpDmyLoKyOJyfKI20tJRnrAAlXabQmS9LKnA
nY3noJ0QCWaZ8cGQYbGbkAIleGseyyIsKvprtul9HzrIPzBvSC1HQAEjrd6AaPK248ACskZT413S
2H04xvGzlqD9I2UY3Ru5F7IQWsLn4wIJERaSAcFV94kq8nGpZYDoNM8DxAPz35g/v6ZPbE7M+9gh
UoMBV2acw4VMp6qShRrcse3UpWtqyMlLhEGBJYSBswyS8epiTi7XE7ASGs+/tl2wPhkLF0ZIF6vv
VaMmhW1LFU23YYjr1JD9nEHUfFirpSBYD9IReuNsWwYg+wpuX+BC+OFdw7uZGEK/63dZozZ4SIeA
xa/HSs/Fpzk9fNawuebzgKDHfQNqm/8AfmtcxxRFd2cpmUhCDtw8K3YdhNYFxQdbHHynisXwVd75
miJfKHdC0VnoVne0ce1g8M4gNP6pZWxb6rebjzQXI0/HNB/WxnbH3UxkChxEnV3tHumHC5dZV5fl
ocbemHlK2lyuXSvEoACYMBtefDbm2c1ww+H3KrWDklTcx4OAWeWVpIrq6ZOqynbSR1thNXrzW+VZ
fboFu1RPuKOTaFKI+ziXQ/Wb+wqIErptKbNG8YmUwvk9/jTh5Ks5o1u2JbNdxruARLSDdCSo4kWK
IemWkt8XLtWswKces/0Tv0UrCMqlJavysAghasYDO9BEh1y7buF5DafDF9SCD+xxhz++785FYfYc
MjRSy6zrGRp7g++8QV6wHbggkLR+7/7XiosRpn3SxtKfbkH0FCDUo8vD/9w8FDKs0tFAM5KI6D65
iJXWKOAayEETAX58GF7rRmwc+wwG+545XX56vtbHSQ6H51QiFWQs/oMNek7FdScw+qrpuubz0uY4
ZQYFvEac5FA9nVgKksv6SZzcU7IUtnf8UwlxL6Ph2XrB/FwTP+oAed4XEPzPZaqVFScb2W47o3G2
dXJS+ZlvmIjwEITPNPc36GP72ZLkwVHrOw+TcjGrLAXcrRP7WKpYiOAgvM8947iRwlZBKPHWyfQv
NllOSRAR9FJT2jQe5UmBoDH4FGOxht/AUndAbG44Wy9NP9Cv/N6PqE1bKn51pIvMq1wH7DPXnObD
Ejm6YDBeeZe8LwJpp7eCgp5Clx00PtXLNgg9wKLTH4f3RFl7giA/dZ2GbRb/UL4MDr0EEO9RglTa
+TcIihVT7krPY1hI5CZg9hd0i+d7CWjnkmN/YRdLmCoDi4BzBfwC/QaGVusbwtldIFc5cRKw8/4l
npRtbdyaqIODEoeEKCEFgoM5OHJUDIVPx/IDYP2FmaVGNq7CSkaG6qXQo4wCoN0HdaPBEO2EB3yr
phDiF1/omVOHr+fow56O95OtsFQaSqLvHst1H83/yA6mO7x6cw67r38IqOdCOJyXUSd6R1sxz4T2
PvyEu8uKhS5/c07Yz1juGhrsiB+c/0DIMZxrz557tG4j2Lz8h8CqslPIQFDR0prXrn57ZSXQ5VCb
F+m2lPa9MFMh5nlfCZ0JbNB6rKrSqWnakjV2G5wRP7yzxDX2usZ3bQXx+iBr2J6wyT8eemwR0M9T
phzhOmkqPquxw3DSJJzyA7KxCLV4Iv1e7OV9Klhov/7ixihq0iJGpe1XSHMdAuzcmFWoUmmNGYkj
RhbGWpd2I9/fe82Cx+CcoOEAwzZooSX2jE5dg6vloi0MPEeeSExeLL/tMwlg8AMpeRUH0YnjpcUK
VtF3MD1aGX5fWsqFqATkFZ2oLjtyoVMuNwllT8k5gAbzheylHrCpLlMBetWSpb7M5itHL6nYGhNs
r7ddr+p1lr6TZ/g0Wbjixj+bMdnMuZo8LhVUilaeEyjtXglVhtCk4i2wPpQ4HkUu2FKVYKGPNev3
Bm5JhS1i+eFE0ARnNgAoTYlrJLXUdowOPL7XwmKpPzSruAw0NzGvynD1RU5FwwBqwuLALhf+qpN1
kbbazyvFKWeoM6/TzOt7OV8CaLwrpfgiuEtSzHLOxKF6VPR1vLyeIZ6u210rVECHEaUiriX9RqYt
mJ2OAVhMf0cBjccjKCvbKxasnCafke8thiyAC9ijvyn6dJYAodWXEBpc2daor95mpbV12KFsjklo
Sq2tLMVIhC3yWytAVtTTTeeAPzDlNTnxN3C09UNWPvbywUd3l7MN9EhEkJQXBJzB6rtv2NNGZ1p7
YIULdU0XvIz/xJjajgN2XGdWTZ4eUcXZVBotg5BmS8B9XFrmy9odW+OsdTyd/j3uQSmzHjQVy7DC
JOzWkyaqZqVVrOxevcMRQkQ6P5b2xPGCEz/R37qklxG/o95T8JwrYpwyBlX9z/z6ZyGY7VM+dIiz
oPbI0qtdizBqfIgUQchOLlnlwEJZqRtm88J+37nLWkugdpoVZyT4NYivtMurh5cN0hG0W495k28b
6vKDPhqx8IiVodGdUb4GxGcxg2j//nCdnk+Gjpt5J0drEgoHZJtkVCkGqKJpDc9DVUfd45W3pa5e
K85+BuVDoFylBr+6EommdhSarSvZ3pKTBK7xmnUIPrpKIkIqTkfegmnp1PgCzosEivWq1Ylce+YR
OdjryP4kI8OCchQhOD9fO3ERxDycAE2cU60G/pP6r79wliXRyOC7nOvbcqnrRwkz0cdIlfGfu2Rv
+CrgsvtwN2Exyf/eOmVBNALobaJ4JIZz67t4DNO7qklfsCMysdM3UeMiQj61hEMicc3bmfIqBjuN
IBLt9L+UecMr6xM7yJloRV155Yf2zGHfmqzSgcwFiBqrntDvkQpMCeH0fmA2xqYpYNXOfzDI2oy8
iFI38/ljdQYV8bHV4p4yvLKtZK8lKEPcBqoUceQ2TTzur+O5y+r72WYdX+MOSKdkMt83w/QOhKZs
LQIbJLrek6zTGMFtUcSNpav8+NN/spj28RxJxUDQUBH0+eCc0fOzHxFtao439Kkdxt5uFK9zzJXW
2vwvAjmJBiiyxGFY0nLt3PdL3mabWfHJ/LYULot4K4KqC3rE6rOlUqP8jRIbnbiHf916spYGqOSV
Uy9DmFmLtEwv3HWeppo8fUU/lRGxkri3J1s+/PEtKIVJtG3D6pMhJX74IiU92phr3V27ld6etzLm
n6trbPDpsyxHS/m1wyYBFI82crKfxJwiftxt89Wh3Az2fsVNnNBY8iaDMQWgVjl2kNNidqttmHEn
Dl+kBK8FHWw/e442DM8MQAItifCT70D1AknaRs3lPRSNFLVjhl2Ny0i+begaRVtHaM8bYTciJO92
tGVx1Pub94vb2TNGc192APHLFjr5qFz9Gbie+k/n27qsqclnrIRlyHF+gzbdE5to3nKJf/7MIi6M
Ia2F4iLnb9aqyNPlfQJ129dMLDfr4oUvOOajia7DBfNi18iNfy9gwsgsyLcpJ6pK5KaYrE55njL3
sk2Q4WLsDaePGvqG9eW7b/mGUSiALqM0+vVYIBgJzXGtK5Cm6JVfmtvxYOYb5iIPIZ6VjiymBIiB
I7A1j0CHSoSxAucAv5ZA2UMm2xO1/RAMrVPgMF5QgyABeeTnIYct79GULPYlfh31wosDkg85zjOD
m7Og4hFiubjMJp+6giLqP6of1KcPtHJwSZjCx+odXCj/mHOboYcofZMX+muEjqSvLhU+5efARM1E
KTplRk+C9Ow2ufS5/cNHqqlqwO738kp1f1AO+dyBei2hJDGMeC8gGoH5yskUhb0so+2ab/OM7/OR
xx1xEb3TLJYK7m4kQISwy8ao2pbk3V3qgWsBFzC2Y5QnceadaintivQ4vIROGbQv6EEQslltGwRK
GL6Z6KR3QF2jiXN19XD5N7/2IxXQXERtUHLhwV0Rua7NQpygok4WwcynICHpyTka+yJZEF6OeJrs
3Ov3djuV5rHf9iTC1zmoyKG6gLSQtLaKWjhElzgOQLaZ4hlUwEjftbaAxUEFUprUnGb7FCggGe2L
QAvXm0tlWhpMeJJAx0cU4mmb3tA57OGEzZb5AlMDFKmOEqdEMde8aWwUHrE/V/0McO5ENpm54p7N
QSLIajhRpcOqhPhO7ZJR33nwJiEccl3fPnuUjX35P5Wt+AF1KC5PEJI7e9l3rbBB8C4TNeltQF0c
eUJIw1dvEnUZT/V1TXCYnrjIZLVnU8WSMOu4AQ7EvcQKf+eyaLthpCiVmzic7qX/zqSAe2Yq2k/9
n20JnMYgG/13iYUk6f76Qhr9i2oA5lAaqIR3cJQU1I90nYPJt7+H/08nC2USK61njKeAK7gjp1As
7xU/GYMmjJaNl7YGtAzDTcJ+/UAZ1cuPqNIEyay2NHYLq6hhyGX/SXS/n0CACofuXv8Ep1dECAIt
mbaMYNZPMJ2Z7+d7PK3v6dIt5h1ah9wPH0rXrSjusjGzZ1N5vLLnhqtqjLsc0mh2Xtic3m0wpLF5
glQkXwThO8KERZVdQgDQ6MfCMejJ8AI1OEqHb55Rdd9eeLYbFqh5UKcd4cwEaKBJmXuSiJwPXKE7
W4YdyYGvPCA6D8ST9Gjd/24zUKhv3YOh/49OxROLLIHlpeeGd2NkDnYV3uo9NMoBNRq3iamnJIku
Uh0us5aLNxc3zbgH5it4WCqNeEmRzqFKc0kF1vrp6Cnq20DcB1WQAI6N2MVcX2vYH0fbxABui+wJ
kM23X1crgEmvMdp4be1OSfro4qMifgP0//fcdi1tW2NtT5gxoT4b6V1Cg7VkSb2wJ2sncr3cu0tO
s0jlFikbiuhtffflQSGC8TcXthKKHgT+7cyFz93vCOZag40UGcYbCZhcEmXfCwQuAMajW9eokPUY
BNzVF4MqR+cOAHwmGvvNDzXA3a31ur3RADUPZYn9V0wnspaSDwZz1jlUekIAZ/zlCyheatUUlNER
+LuYGdSyIR/3TNjJwwtH/INd2k2nmrFOUIVwaovFxRxqzz2n7IpZYo1wOqOgQnyHqLI+LWilZuAi
TMMZz3KxjYvip/6gbFL42MGrML+23ctPNcpxsv/MaUSitwiDJkqz01R92NfzljRCaRvE33y4fVWI
8XY3ojjq82XjcfMTGLhuVfI/KsWg8XLaOZqWG5Fq7VxkVl+6r9TBQEC4TzdZl5D6t4dbb+X/zuC9
NNnxArPha5oD1h+7ujxZ0fTPlU7UbuTbVGcX/DKUGB4yrcdn2EQnLJZ5wgD9A1tMgQlf7X/cXQFP
nR+sVTg54pByBf8q1K1y5Ijn2ZJSdx69waqvY4Ekb3foLMgQ5xV9EupaU97QZx61a2HUm1KTWo1t
NrzVxidQhnHSYH5g0S+dDgaE75M0/hv065c3mCjxRYvcEcXsVB4calZVUNne5v+5umTjaAdLH/KX
fgL6fthC1nUYRg5Lnwlr8AO68SuSFbJqG1aqqQKzm3q7LGBQITTdXlgQRXDjiYO/OxlJAR9Aa64h
8TiVlVAO8Tzue14gmSvf3t6QOQogDD6yh3914yvEvGKCzDAoeRMvcIuWIpNc2HqqLYSUbFZrg90g
eRJVyexM20J7oJ64LPEsI6c6+fRatKWLVvMFGCXB2zJ6eQF5IYbAu7PZhVNksiSiyBzZmVkTSrMS
iziZaaPIPAm23zK46Fo8S09WR6W9/g3+j1t8vHp3/mAoOa32+zC1nD9veuGI9wxEG4p/UKYQijcP
W6QLxWOmNRg8m/M571lt15ePUQNTCJ4+6LPrV+OwQaiYv7wtXVidlZrjHJ9D8qxUMVtzuR+xeIsc
pye9I0sSI7eYnnuGvvBl/YmR+FQ4Ewkuifv1ABLsnwKSQYoPo5tR1p0U47JAsj272uVd+nelZs4j
tWiQEoa9gmOgGF0IXL45Y1t7Ez6Sbd0kBpnMF1+EhimS4FGkm9oMMkrb1HDnXJNmFiAqYBofS8i1
kP6nGeZYj6Rd9HcXvsabVuXAEJoofKCzqU4k+8E3XrxY9A0JYsXLyjE477CwKPh5rFLm2CVYM7wh
hvh7S9mc7ppYjCcPUtlhXKkJ3Fa2AMyFzkiO4KMipxJbnt0ARYwoKOkA9N3SPAcfFakrPpMU9II4
3Iq0ue+Dysqy+hO+gyhR0ZxcHHzYCBA/Ei3fY1rwUH2R7Q7XBWDPXzIK0vLVieXyjsWDT4TLabTe
/kBT/YptNK7aGZSScxqtgOk3P1Vhgx8NNu9b7D54PTn718mbqwGMzFE0mlNoefISiVRy803rQoCH
hpENKtQEKXBaYtBhKIb6kx0C8xyqESdMfABI4KjUGcP/sIQUhzeQztmsVveaozdw/24DGBKSgZQ1
i+SmYzTtvLCWpB93UvHilIokSpQa8eYslU1sJIiMwutCICdAh0esGLDVHAhz3e9vgzfaqxIU9URa
Rh84ZTsZrgYftHl22ivlAuQWBIEp8xLGjKwpKLhhdaSWdLTXYnGcEZ4vAP+pVRiWAChPsS+NPYuq
qGWbdK+TvBZQ5VzuCzEVK1okUHHAvpIE+dI6uqbc7E8Qmg5AUksnGjANrB0YSGesUxW+4RxqVSx0
BDmmTWYpgOx+8PfKwS9p8UpevHK2BoKryD77tJEVTxF0d+MZGLyFSp/tMhtyWnyj2oA2jZJ89+43
o0Sznw+sUpgGfd347c+/8RJlGRIGRBOUuCvvcppkpK+HFvakMhlx7cs5Kkwt/gQodsi6k8XGNmE6
33k1lviA7aQczsXbOzOriK4Twk7S2EsEUzznjLTCTwubDhMFcztsC1zwm1kald4zNnBrPKkPGV5V
gRe2T6kgKtWqdK3W+FB0Ki7zn+oZP5HmatObA+AjZWTbAAw94JJFvShuNRyTqhUt3VTIrzA00Sri
wRIjE9qD8yU1gFOwCCGI78FMY1+5o87/5Dkw4KBe5GE/hmOP/CcmC/1DW6Fv7e2fuUF+hzc5w7Xd
ZNfTkGfvbfX7zwsMHmx2X/Fm20i28MZnGFBJpeHEzEQ4oASBWD22jjxB24lFZYPFYJ1XKHcmQEeb
0GjU8F7OvAhaCm7Ky2LX5+LyIn9ohq2m5hbLqxNuwEYE6lPmc+3NcIAlGcL8yg0ibjHa08/Iw/e3
SSzIO5OsPsbNCGwtxik4U7/lt9wieZNt03+2/l7k1ZSu3YmRBMMC5TsUj5Ok3U9iQUYZ8Fn2zlTw
GJLM3eOhnIgs+YStBtgZTKQ9ZKhuTwCYV0+IEWLeQEnTF4mQmHW0ZpFgZ2n7wCWmDCdySLwbFQlN
Hgop8YFcT0fvp8+glsAE/q67euOyMTIE0eOOAiU2m5r/EfaS2nCq3IqFJfjlW7dzEuc2OMLg8Wwc
QLFSwJF5gWEDvdAZ15662k4Z2+DFNaxd1hSl0GKmMsAYTL6rkyvKQ7s4jZWyQ/brcJ/45CmVs/Zl
Rdk9OJ2/5YiBDn5sff1sUMQ7r72cYOO9/qWHmhFmDok4Okb8mN32VOFfg+q73b1QQivnKibqYjG4
JVuvyFRm+lPaX6FLVhgTdoL90svIFmvf6phUveTB+2piMJ0Xs6JIJ9PcI5AwTl1cK2vIX6YAegeI
T1yPA8FDHrfa4HemPtlGz0fjPuRG2OQiAf8ATvILGODywYoQmZ664deTjWcwPF5FsivTCvNFgVRo
Wakt+W0xBrIWXdwhA4Y+dlkB0iDQZGpQf1vDyPZ8RAJcCB9OFWl5tx/u6CHCLHGAofnPmNN9q0Oj
4n3C1sX6u2YetNA02MvQwghTmJRYAH9x+888HCzcBSmu4Gwaa6s+k+jNZlqtJzrnpXAOru19ePT8
OhCTROroq6J3sThvTgyJs3dpGp0HZIGyjEkHTvg/dF+mQj75WyD7Oyqeg6y0lSzG7YuEhalDDDh5
KPoLhCm10AK/8mNz7sP+fXxygeKe5SUu7h/QpZepX0C2D4vQQO3+6WAwU+UHIC1SL9AzP9Ajes1X
i/41V/3dEgClzRqEiHn7ppVOyLPFwPP8ODAPnfIjSQHOU+wQ+snYzHJjXnZnNbroQm/RUtwjwNcI
fjoecciUYybrBPQfyk7vm0QQbyyOk6TXrgPTw6rpAZy3nWLMoc3U6AMFrqFFgElXf21BaOCOwVPr
MS6j
`protect end_protected
