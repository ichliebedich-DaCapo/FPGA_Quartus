-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kH1RK5LZ6/nEBWGACiH66+U+NHDAeshtRgKrLMNB8JGQE/J/vqjYLpjB199OOxNvUQa+jGXLavVK
D79LeSgpNgGS+K6YX4GyytiIMjE6fHZfy/QAxte22Od+6dHVCvzxGe2GTVmCYvOOOz/JETJAyKIY
AJ05LN8giahBIz1fdhcypNEmVzNJJN07IlKi25hrkgqWFuzmIcEXqQDoe+qcW2zJ4aH4OZg7c2Qz
t/H3rqL37K+iMiCtRnM5mEImu/+ZdaalXPvjNR1Xfg5RIrBScOnsWG3mwJbQqpM8SeYbaGZj2+DB
ljDJDiKEBCyHV6YrpiAZK27SWuh4tmU7gDQwaA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20240)
`protect data_block
JlSTFJps1UJqguqZpD4JgCgcuSJWYo30NyMkk3gTCGPDjn/B1lKZW/e15qrNBkIx1xnsRHGPflTh
WOYziahgyGvqpg/a2Flz6kTvD+A5EJsjD1nrBFKt5ZzDW8NKaEr+sWoH7obYL3MxRVPDT8KjPmA2
QZ1HFvXMpBWVtOAzUWq92OxAwe39CoqRVLB6fm4pQVxVRQeXqJvNYJXefMq0R6zg5hvT1S6dG0IA
mEbLwxeS9khXuxsOGgECA/7tgLl/r9ijPQrzT4ILUQRh3YlKLZ757ZuZvZaDigOJDkdHB21ZdGcL
VX+etVV+lhUIvDhUipKexLSWEJJYF8ofqiskgEZh1ZcdzUyOHd9+0Tc+ok3Lc/SnaiLtdrg4ylSg
eq7ebJU3phbcupoJRTKiWsZMh3Q4Kip55723s0Gui9atcgVU1YAsgjD3+pDG7CVBhAkbJDhuX/AL
z4HZQRlErP/+fKR+NMW+/HRv8mC2W3UqWp89PFgwwC7Ez1qoXPk8gMZceEfnvitCXfnZnX5inuZX
dnZBXcpwnVzh8n9p6QTM34/Ieu5+aWPx5gejs+fTkakSTwpf7QFG6+o41oOe/blw6tBOaWFGyImE
NMkynXJYAz7we6CZNbop4c6kDyQGrtTjzbBPzQDR1JAIZJXbbigffhc6XECJKROWl0p5ShKo6DoD
R9G2GgePrmArgN3lwcrxIQwmOVK7MQAfB8ZwZXf34q7is8bHl706bJ+l14Gtf8yWgK4CXEkMs63m
pi0OnwjzlpPGjPOLKfk6TAR7R6NvDBCHyOq/gJbbmoZ+qp8HtTTPfhHA4GfhaVid/SHH/pKuDy1t
ZLJBrkttdY9WeuuNzDbnDFV5hlCtxxB8TOe4K61KoxeSvDvpkLNwdXOTdJBb6k+lMKMvpSh7h3CV
iYPnxqfj9mr4mt2qdoBUhvFzOqNFwrT7t934U6yeDVjgZmh61wbeIz9Gtn9mxfXuS0NagsACmyUJ
UbGxX/TRy1FKLH8FKkQyYPwUREKgtQBk70Ri+vl0FEPRo1UjnlAS0jbbfR0RSeX23J7xrLfkG/38
EibwImKnoHJdBOjsFK1YaeWmEoSu3jCrPTebFHkhuRNEIQOW6ncGdeF4wiIfeWTkGJ66FhwHsjXN
LQXcscKIuCuh9eOaV1AQf1VKJRjgTHQfb+G7Rhfvx70X4q8lCkuhe2yzurrHc33Y72iiVn9/JnDO
1Eruukm0WjrhEVH8aOUxVTKcDG+kMcNz3YYjMHsNIxiyIxm5NuHK06bcfCQqvhvCh1IxG7THaigS
wmgGITJEq81DEkuAY6VzlkaYHFXsAy61AVkyC/YEaZBVFsIB75yAqVhZN86AeMy1YroKmfEmO8Ys
mM/Rhfo2G0vfpRYAmLboeA9A4g10HjWZdnn2+IZl5Wdn729qZCeK10EAvbl/VBF8iXcV83VStwQg
JHNnpW+9FOby+utKuuAaqmOVKNjNqqEOxAM3Sxly7XNwXBmmd633lcz5Wtc870DaRtyBHurxSE1T
EhSb3ct1v4dVJJ/CMQxtTbuNk3GHrw1OfbTcsY7eF0g9YSArQgslO5OPjJzE32lrUFOTI8Gmrh2M
KuAupZ0bMDz2eGEWxr6OD3jgnZ/mnwoMw/yINjk1ZbHIMp7297wZr8BNIUvMJ7CD+ogXyoELtBph
+2iMgrupD/qG7v5iuR5p8KW5Oc9RZlGKsPw/wLTidaWvzzVrocEtvw+4TMEUsoIH+lkoGrTBT0s8
u48tpocfi7IrJVSnj5D7eWMInrd+YUw8B8MFRuXbAxscn6hCrNXUKUpK9+eQfxQkQayV9VhhYFX1
gQyFP2KYsRxdqY5ekEQkQGnmx+uIvY8T9FFHmKkyTf54zqASp5yQ9aP5H1UQG22BmDvCFpklGm0N
rZOrsx1Z9V3gpAe/DE95iX/eWyuuLHveC7NSYvlguNEgSUOQ0ZdIB6VgUY68cq8cLzwxP52vsMRf
v3ar4Ro9cnfO5Dx4//Sp5gSrxb35ojDixye8I6VFDa77usHprfzfQvSnDoNu14FoLQew/2v11soF
5A5VOQxcrDQqo9n66qUoQzb/O2Tr461DBIYj42Jrc+His0Qztd+3t+wk590csQbsjpqL7qwKei/k
X62XRfwM/rcwqddIMUkVz5a/5hO5HGhGhx9ZrjcbOJDjHljUoaJOZOwN198lIQw8Vphijk+T5qj9
GStcQq8ZGGOTXGRnZMGdulO8AeJWAJAji2nCXnbQ9bCNNHj4kSl6qYDOnLnT1Nc3aWn5pQAxqrQN
4FxarzKgb/JWEJmMIz+jWgUhgma4fjjPthAYq6Uvn0XWfX8OWMSCZ54Usyc/1H8DRIpOnwFGX7PF
tlIAj8cIn9WIS62egzFFlTUsDWIpskBsmA7gYtD1QfHa7fx4xtRli9vRtWxnHMuJy2yesTFiKMxw
tlkT9pNtzRW1lnE6K83aapZYnUvtAWvbVfh0oV/+v7vneMg6LEHWaqLlCLdtG2r9cpr6YsnS9/+J
suvvsREmlCb9reGBhe5wvSYUaz9BzD+NIgnufrCQcuXzOfm75ahg5LsCskuR6qUrHLsYd24I0VNf
urfQ90eAcFIWFD3JLbNowz2d8zhmrtZJVfF8kUAF9eZbywVliMhzXkvHbpfIOBreIMVxvj8rY22d
Ye1oaEtCn7gUxp6aK0JAu3pHIyLgC+OyHe05BnEFn5vx5sMRpiRgvRyNJwXtCdsmxjyaB3KhFNLA
anFvOtkK10mrZTjc1n3n7xCZKg1yMxwm0uRfRw4s1uJkZ8lbmYD0vBO3skW2ZY2xyRsR9jUUV7Pw
Tjtt6te6T2znWgjDTJ/WatMc/fAXNin9wbu1msl8QvZ8OkuriPljJ5oyypK9azjLt0hBRvZRIwxv
D78fTwin1dwiHEjJaROr0Vw9ZZwUHI84883BkMrcsh5CBbqhjBEvhsqjfHUo1gzXtRUq8mkBFuQz
SPsARJ+5DVJjrSSTdstrfy5Uae9XcGA/8YUziHjHJIAq4xx86zoTMWKcX4WcjSdRyb0SKn+5JEhi
GbbWodrxdlAO8sllSyMGwahQw5C9sK5ByPc2RHcTEqm3IVa6sLHr0mQb96nIzBJUfNecVcPUVM15
Bt8dl9dlqWYhKp06dXMezOOf7jYYRHybYBMHGK3jfMFFQmVzqzMlCnUzvNxrXVHFy9M7qQtplNSY
Lqa7mkkCXv2/Z5pEHnbUYHnEKPjlFZUOGHDHPjH3RigjH5wBcNtiz5yums3vY43GXZ2tMCu4Vdo0
7/vh/VuKKz5Z//91dQh9P558aou/GcLrKfbfo1IuoJ9Xoz6CHDcpbDO6O0AlwTtNF9A1286HTBNx
B8lJn6ylUk8OIMZP07sgHznrSAVqUy9/JlEkxwPxOLxpydZV2PxsaI/5hR4HoKsJd6NChI7A71IE
ON1gtMQl7DpK4x6xxfxu0zlRlZ82RYWXwfSo4OOD+JQH2zijfIg0mo3gmag65Ch4mKL2e/CpYtaS
BU/hMlqFwOWS4eS4iD1FjsjwlBaopL9UqTGpb1VIQ4bBkdzcIDt3q4FkgthjNStb4S6pFGKyXLPQ
qsALlDqxynl3uOrw9gOIjF//TP1gtvq/aJABUCxupc3EqXuNw/XRPK2OKdZ7PKXHfTL9bAedc9ty
sRzYJ3pzTTsavOygEeMtTUuIByAQqWreGF/SjMZi66vjd5KY2xBjzZ1DsJ9n7kxT8798JM4r1i3m
9LQz4dFh6rm3UG54TM70lrBrPOdQp1eY3OoLg+rYilq8jlOxwpbXjYpY9DJmv+y1cL2RYRrCGwjx
HrzSzg/XOtqSjPu4ZdWZx7kbX2BFrvoJRHM5AJnM1NlJJzQ9uREeFbkNPA58hGKXBVNdWP2+i8oM
iJrW47+ONKEcM/qGKqF1ljiU0c/IjqyXK0fftnEG5RpRe0Y8kmxqCSvO3vm9FBh2e9+tgH27sRYO
4sno4sN55wtDIg0lU3JspOtkstV8v5nLuFolfLfAt0HM+p4SHZ3TWiStMIUjFxr82L0tPY8MZ0W2
jFgZ+Kn83Wf7NzYHo3gqHAh3XYsK56NUZ0L4DDfjjhzJ83g6wCOeYmF2m/pt4OGf/d4b48MPSD9p
4X6sGhtiYZ6ZAD7UJxpuhRUuqRTHJuKeo8uItqbHLq3Ty/hlQQ8iNU6mRILMlz8yMiJewB9QXfxF
0ZXdzfhw/Y44GNs/UgnOJJ6ggsuuORdgZS3bxbksKhCpaTdFPTm0aBvUTUt84fro21dzBBqtpw1d
jR2oRgBN3YNU4NSBCRaxX4xfYSC+SIKiH2vvkyoZI16240XbAGUpJqpQERq2B8DMD5CZRvSVQHIF
2JktzppN4jLzsIcS3JM3qNtsyJ6n7ySdZGHtvuhAtulZCqNy3YmWbd0HIVf+JZsJslEJ7kQt46cc
LhjXfiGDBVAway2qBL3O/r3u5gEYofv4lVJ7Bb2StyGdbbXu6+IHE4hwLthRtuP/IeJep1u8sapH
A6cmp6k5SeumZYvCRXnMqeHPQGYLrKykRd3DHXkN2UVCSPp/tH0xZQcGwnVun/4LGS9uy7sRZdcB
U1CmruVfjdH0fZaSVVvsGI8xBNKIjMH8XFWr/jJmAGa7I7LqnIAV0X8RtV6IheADD884zXaMFoIz
6OCgZfEoIE1K/Qv8lqgog0ucJxPxzR9i0nFfkmi59tTKw/u49j7bzzN9Lw5q3RCxXjr8c1ATaeDF
aL8K9uOaG1/vwO6QDkkfk/7tTPWePwnRcrq2QTFxmN+RlSJI29eMiGVxb+P1QiPtMogmII0Gm/WE
02aQ/qk/fEG2jG3WF8svGgPx7cmFTyav6y61tI+bAPCJnxWGBCw0apg4BfO3sw5v4nNP2oBNmodg
68eI6YlB9I/rFRK304LyaKbnYicuqxkEdjd2N70jN2eRfSqbNKuANI3RXeKk0AbfDxxDOTA2aD7X
Ah0PcFBjIl7CvDUVAWYB3lldj1cu0PE45v25umnI0LbqFTRZICrJbP4FEwiKFKKVYZ7hEPTKlm9C
80rUNUVkHX1GluAUNy8A0ZAwW8W4Lfk0h8HZd1WhR0OkRjFycxY1XW/Otp5Qs4aKKJEEP748iQXL
LrcspL6phFHBQla5LKu2dwwiiLlEj/9zCtnrqunejkg6F7LbVlEcHVjI1i9u3UCz10x7tZR4hx8z
WXh1kly6PsEqImVsmXZjS0sPKNltI1+ScyfGBnu5gKhsHrvYIC4O+rxRZGajKg36p8sLLq7dfk9+
EEgKoD9vJ+ClBdSi/sXFSYzGhHLkLFvSicC6F+ItaL5X5LjqhPEMDMYD4Z94btUVAYBdlMyeIxij
A7Za4oJkO4B+3XJngSwkiOaHeJGb2SV45TC829Bq95H4e4XEOWwSeyKmBSN4vgXMefThmn9kZHZJ
1jAszczqTqGYdjwWLQPx1JM0a6O5M3kHoGIxFBH4AcVsLCJ/ZyM6KJzhljRI0b1A6VM2HbCifLZo
/VOK3v1nm8y+2hKPV0fVcDo2D1ONKDMB54o9BiB282rmK5ikQAXktO74e+fYV2aqNyR2Y1hbaXz/
fz0elGtWOXudSB1hhJhXyjw0ekBvbBsuZb7BcJPFJTr0z5M4UROYieI7Du9tGxIxRI052t7HP9HL
Z7Bk0PmdM6jH812jAOp9+m/vItbzv+K4QPgotpovEgL7UygRpgRU2XDZpO2AGnQAInq+zRSPE6P0
sj9D74CJwEc+K4U43kf23vpD9jLkQh8jaFQGPQurX1S21GuJjP86qimpiU9bJIeR49Ul/3CNdWjU
IcjApdyhuvmnQSyloGSd5mVigNdSEGJWknX9lX2ZEUJInI2wZ6X9kZ+2y8PORCWl0jaK/sVGY/UW
2Ddmcjeo0KaVcLvORSP7zaakm3zZUBSZaVSgoIKSNM5em+7Ce/KtyCDn8vPpOzUuxSzg980LEZMw
0kEZ5nSlx1pcHjk1s10jy7DJGg8oosDXhqLSUg9lN6/2fY74WZtRFvEt8Md2zNuCEROepNe3b9ow
IAvDRj6WSnwxAuybK9Xn7A630QNvRV+AKE+QN1D526Mb+UiEgaN3IPRD5oMft8CMEQY2DenjJzfc
bPJDGPlybLBBP3TX2qT/ZSCVKjIaNrNPVC2OrVShX4FkrUqaKX9NUlUcvrZrqtgLZLiLlf82xAsx
UerAvaWqpVsxKExRp+ZrVtCXrL9DMA7RI00VpsDffOgkg4EQCl87IbAqDupQSD7cgnXwcTOGlkFs
ey/KP0/uUg3mIC4EUIJLaJX7clBhbLKTF7HM2ZkRupMurxB37vUPrLybQpX3Wux63c2OTjMnhke7
llxok39XFkMuZdlvA1t7utcP/JcBrtJI5W4uuv5vxYR48pB1jVvpYEL8AIIT97JG4jn7P1E+tHEx
ZFnMNMp3+SdGhjU3azl2H/ZZ8M6CjL3BW+K7leRU2tpHf9Sqq8Dll6EF7dYhx2fJtsUpB7xuGDHF
ZNCb5Tb/e1vRg9G0na9xHEGuRFfck/qvwnTosL0dVk1gz5blt/Zs6gQ6fCmETsJLSxaFUhSITy/7
YAlJ078ANiX+urRu5fDL6v+5spcNOZFrys7w5KFItFndh4qDKrh/Bij3iswgTiwSUfyjbkzSYtWi
bxEwlcB5cWbPEqrhjIGVeX+whXM6Rw77uX8c9A/hRt47litZNXSC/VsxSiDYa9xjATqotNSQB2E3
fg9Z8AR65cu1v3Fi23nkKHp5EpkDeyL4Z+5+p4IokfzAnhhqtCrl/0Fdim+mTn/pys2zCohtN11p
BVHWa6phaCucuEHletcJ1jA2a5jNSCA94oRquV7E5OL9Ny6vfeVCK/8F+sPKgfX1ItEdntfs5fgg
3qAC9V4OXhW8peQc+/4O6Ye73ZhZbo6BgkUxieHWtTDNGTxEWFj8jEMP4A2TYNjE3JxGg7nHapO9
zeZCmimH0M4Zx/Go45QvYaz+gvUJjez2nnow6UcrjLY33M+kdSeWp/TqjQ7DpAW74h6LVQVwO9kP
yotnUdzbDYySqA5W555zBwt3yggxmY/R6n5T3A6PQxEZ64Qe087XFCgMPZNOrd7qJ+tLfGEqSa4D
xfBlvaEMhTPvbCmNIY+1eBlFMygb7/nf5oGKr8ZfSCqtqURXBglCz9ntl9P+LrTwovPiQqbiYePr
nimRlpDpVaGqSO/wG1m575hz/L62uy9Hfc10SDeV2qIVmvzxDPUFKvV5zUeMoA/6UjuNl+MALAxu
9p7FZipEFmywcwu+apzh0CjKNzBLoeaKvDK6CGkxC1XMgBh/K33/cWbCPaPKtp4sGQUc1V1wvJwB
a45o0kSQIbqWSnt20lzLe0/WesSmCHX58i2zT7toB4CVVH02Z0wi5R4SvgauxjSktf+ZdyPdh66v
qOZpElGWjGPIO/RbxZfv2kfVZIgV+XeOKYYzs8OAQpwbeS3FIopuXH/yHKwJfN4lR7vkat8bMvLK
yF0mxVqG7Dpksp9e+4hpythyPxMj4hIZ5TbZcQtaHbdamHuIjDkfppfbg0eW7wA6jUJLFvFNuA3o
dUrLseklIcPs6X9kLiWM6BPgUC89sQYOfBFpNTxzSUa4ngxRdS18L/n9fs3jV0McEqRL4VhGGXfV
nLIUOjS7DHNhaeJsSJwMN+R7y2kkExyy2wTVf8C+B2vXlBDlTnsZTpJpioPW90duYv1gk6AwDY1O
wnxvdlZU0vGc2sLLLfztFggbxA2ljMmDeOAZcelkIRFq1404nom0dCUPTtnftYlqPf9CbdqNqbuk
3222Hq+avBoPeObVNuX2VLVVJWYHXIwFYxWYob9oYuaNDl6FYMZbRHK3+P1HC8o3N9mQD0jQxZJ3
kj5xxBnJnJJ/q8YXS5pK7vbmHpFSeBg1TffCDi4XUI0hlSC7Y8EoEzJfehkJ/0tlnH5JYLVNT+Xv
ZntzazkBAhs4zUm8lBsMkTL8aRlgTh/xzepXRVecY4cMDuZ0gUahKFtu2/07EL9v52pBV+Ce6MBq
FcHk41JdnEjVtZrgucmFW9QBRZmEdCMVhb1ubXijnzyODpiRCuxTSEjC1bW9G3jfpcNLfM4nuXe+
2mgyCUtaUPvO8phF8hIjxOhTcXisHjImCU0YoGc/8aJcPvF7mdm4A+KtnZlRUzlHMEhBAl8mqPAI
bkQIaYmHaw22L88e/86jw9V/h1CFhZbhbZ1kraDUST2/sOCYHgXufQn7vR1LmRjqdBjTYbgQATab
XNKfYaDTn4WdAlN9xsx4xCT1jJC40UvXq6gVFWR/9hpfkyMn/wE30MrJgGZ/zDK86ULWJ6+1TUMO
ONEod7NkH7stfBhUku6NX8HY+I3KbO8dVKiXtW7q1o4OccEDBkr16k4lluWnxpufquqiKeiHKKWH
clS+iQkT0FIjQs6Y9Mbni41qlkoi2NMBb8a4BO9C4XOl5/rrljdTTs/QHYEGfHPgw/P2FgfGfKlJ
L7LJesUWk6sTeX68rq7EQLDLAbLK8YQhj+y0AlR4jGUccbaL7XG6EHyjlTVIiZp4pPmd65lV/UXQ
htQWaDrS2MynC0B5PnNN46GV0DcyGr+QSI0g2RN1LWgSukL5EcHoEaoXh7aXEpcJSCpmJNcG6IE8
mp+Os9ShAd26LZgIgnxgRJRGya5Lwibz3J1eKbhSvy6UcBOTfCS1W0pkjhxZa07F9MizYONBlBHF
aWWge4NkCMnu53lACQ2l4lCpM1atxak/RfFYbk0nJNGmTeh9A2jOM7ovnsshgDuYboRa0PWkwcnc
wZnWiGNZ4rxA/7oJ6jrDKBukQgf/+ARTp2Z4tArKazAV8BD01FIPlgYbgDBdaz3qPGr252tlZzT5
8GVPyGR78mfpXy8QPM+1QfgmR/yttIyXCAEayXcRX4Bcj3PoWXf29THVgfytCAO15Y3MnhK0dPlZ
9yl1dkuxbTMIoL90ThHu37jYx4U4GclRswxfdCgI85iJZ8m30ahJh1irbzbKQyreGi1IWRGPden3
7nzYw4lLc7sVVJjQ/5J1thnRNCw+Bla4dZve3MeYp/MNbxzNPpw4MAtWcqBzha5qVyIZ96kmsii9
Lm98IqgqL82V3F/YW31bl2GIQODXIrbtRc71ekBNy3zkV9489U9kzjxBw1Qm+vQc0vJMsfDsBzW+
kFiW2YpKBu/D8tmdCGjLGDmEpXNadmo2NHeRprokFqpIPWwdyFZMZal0068L0vfTnKdd7ebdgfgg
KOA0ld0Sc7iIsJunyuEltxLsGcAdBMgcIGCSNVvyda+srkrm+C6AMxw/AbGfwruPpdmF69PYxeMO
gAC4QNGRviUIcVrmw7JwiFCipLE/KMzMHWQPI6OMq322W/ClUE3ArtCp1m7+eivcINVkBXwPxs+7
y/f6EbZKqoPI7BnQFtN1Icpq+vyrKRgiAeXFNqq7/U6wJgfxXOlO/Ajue9O6aVcdWvlSPLrG4YO0
QiqP2QlGt0hZds9wddqxz89ZVLmEw8d8flFx50oEcNUbNZXkia4gicsXDOAC3qX6twkn2dftlcKE
cJnUU5LhztSVir2TDsH+y/vETFDPaDju/5uL66W2ZdZkUzxtg/RgKFitZv9vYc3NT694ypqPnTLP
kfWTeUNb37OZSe2zZhcqjIQB8VBQbl65AAq9VsnrEt4jiiAl3bi8OFXrhcsYG0f53oC0IQZ5kF7z
vLOsrREsQNxAseEcwidAXRm+AszGhtA4pNSUecFhWog/uO7xt4s1yW962Ly3e4O5LXdleTHo/UYP
syDHDJzhoFKq8n2rH7kTqNJAouOUDHeX/ctG0YBxEH/xVb/WrUZj3YpVRkWzpPzzxjrhwuFC9cgt
J+vjSxo5lzkPLvbrdRnqxuHe9RLI+sWa9UTvJpuzDGDrZBsb6RQ3a7Hm7fxMCaehrv/+b28CSlzS
Zi7Oj8McztR6wNGucHqBvssx8s9LARWt6t0PWclbIV0xAsDnnSkfRD+oHqjv7eAnQgPqdg6nzNXM
MlItAOi8Yw3DGaRPnHbImzRHbAC0ONSkxg7AN8Jb80vbsKKaNmIi5ENgxGtpXWYPcIPUBXxro0DO
f0n7oHXA7nPvwa4tb1Iyq05dxJb3qEfSlLSsHDgQIMWUXRtYV2lsLmYxHImObjxXv6YLOYEDFxrR
CiT9SI0vnpjFv82euldzJgYf9J1+xXWVLHEeLEseKrK8OwkxHE55CejUJIpoFRMfD1J7BSOwIcT0
Ui6rDRqcHvFwuWlMmchwSOJlUlEyD1nfU2BVQL3WnsFfDYsKvD4wgnrLyfe2ht0e8F8L3fwBcpVK
xQivQFqv4QIVMtGSdjBcgC38+f7Xh9qFJpAiuPmRJc7qovXizlw5dvtbP7CjeQHH+UZ3wgVJcVvB
pokSVbphAWl1wXbpecRW06r1K4OCFsxxGSZLAv++cVz1IGHEs1ACa9Z5QbFQKUlhs1b0rsWMnvzW
jyhA66liSq1gglbnm9opJjIUd1EPnYhWT8oPFpjgPO9uAoqs/E/8tJWM5/toCc051tr6Opeh8wkG
cxbqoARRi6tz/1ZAyPdDfnObBxHDutbY9nRUTh8JJ+1n7oxit/wxXys7qrXKCtpNc+rf/Lpq5tZ0
GRy3FeQYbUEj58ZmOWy5UEarfFYOLOohmYCP4aeKJ+3xFshG/zpt1leiafeQvTRQiIqNZBd1D1SJ
9U+s7fkQuQudUhcK3NvJ1dxp5ItBvE/A0+LflnspKIObkebElInym8B8NElYA0GRNTIt40diNzTq
EbZ6+o55jopr5wRoYL8z86Ftnpgc5VGmBdnDaDdOaWIngvVszQ8b4C7+dqqs7MiUsT236obLliZF
aCD7iGo85SqgG/4sQYLGzTwjlglPV3lePj8FIVgcJ9alcPdvBGDZqWyuSXOg2JAyR0X5pEMV2jHV
TJyDh6E0yB7HQBMJL59h/cZSB2IhPppuMUoH+orFD+NYGOd9gfSpkIFaskjO7qV6mqk+YrD/TpOF
MW8AEWZuYOdqgBXp9Z54LxBmdjLQoBp6jfEzj3+f57NPE6TZQl51pQsrPn94jfM9cYUGeBWFksfO
1mkuAV6kkVe3Iwy1jqBkkOqrcUgeicD8rUWRN6MJp2wkVXAF5afj0YVBPSN2nMo7s0Cbz+qxZEVJ
vW9F5XbGGcgR5+0VRYHvOCjYnv7f0Z8sWilNx16j0/KRBb5uXVAw/BZPiSosWXRcWcKUDiKJsXkO
gZO+93v4qUiXiXaqPFvAmNUuW9rEEKtU3tcyCz96n5swSyiBFgLZEJZ8Fjyp7pNbQGxAq9XtrUiH
vr9cXwhY3SWMSsA8BnLlJI3wk1lBDk+HvP7hpP9iB4L+k32JQayRNGXMnfZx948LqGUE1LqSUXrR
de+ytMglnAwI+TSr2JvEacqZRhEG9spt1UTT4RiH3UY13OabYSTnIC1EJrBZDRJfK0ST2w9qk7LW
z/QEpKKLX6ijhgyW5RECs9AIJPTBcUYU68WzDMf2Mo7NR/hRSVPOgvJQIWLIVpZFWfXqovvQWejb
hXdHs5rGSAZSxCFsrKuoHOQPo0QuF0csaOKig05I7c1D1tdYl7IdZphudDwUQDVjeXKeBSLfFz/I
1vDr2r2nIRhIrTebKvFLhPHj2wmWKpBCYTyyA6yTcFXnHxXQGdZezmD6qCE/hjprdM1iSg/oS8up
0cAwsIksmYuNwd6e280kr6/An+42+kBr2ON1jcZsGRBLFKipchsD5TRaHJqnDoicZJutLNHVepRJ
bA0ueCuYxoG0IlTXwi2IMglpvCO3cggy/9se87fY9V6ZaAGFDbEBN+9DvvxZ17SduRc69f7V/crc
1EPKb0o8U7tGFV1ckom9uXXDMw+20XLaGsylrP91cpsTcZ6m1Ffp4uqxAVpYl/2BWW/xekUXwssJ
4vWoa72xHLIsx/VrBvtF+Qr4ONL1a6oBXgN0LENFiUrlRI3vsRsNjGzdpDDL6rNo0ae3ry1Sc8Hn
RLNxxzQhD8CvjCAICfjhB4w17N1hIjGRNVt7AG0Z5MXTxwxLTyHrRFd/19ogdwY683Y2IgZSNHvp
WV0+MmttrSvfVMda2b1iQk0+7oStngM5Iq+zGh5xuIcZ0aPpI9P7UeHYsix5v7D8Gq7SZOMbOuES
CcVTsFABJSpUo2FeCoIJ00zYsxOh+feTtc3bJmchlh8SNWTWl1qy99tiHMbEuzBRop7+z/13U0Jf
e9LZmef/sfVi+DdFfdXPCiI21XBfwzxcx0AXlbh+0RKXxBnoDWz5oEbZD7zTArBGhbKxWLyhDaKK
bQFymswlGiB87U9222j0egTcjs7NBmniqIkXjKE8SchN4HfkVpD2jAbzpr18CP9U2x5KN/PayHxH
yQcH7lMi8AldR2WjE1QG/xycY9W/n4nn19nP9aQlhbPG0dfa+o9FlyxCyyyDxeS6rGJP80IingE/
QSzRt7/MY3AGj5E3e2CVpYM3JmPg09801OR1HfrOdQLkHTfiLzpR6TCXXHkxc8w1WdiFvugLr/My
x+huSlEhz6wczWIQ5zEQ4ozePiVteyibH043VDJQB6BO++xg/bfJkqXtjcHNeXsqxEq8T9DaTywk
UMqsuPTEdxzPbDfFvg/WE9UESPVpE2umiBxluYOfGQh1Sum1h7TYOQI688kcXOicIP8ampSR2Tmj
OTQyLVyRaSR5X9T5K1bV80BcZNCdeURYUc/TgvQhFsn6yM16etgKziYA3b6UgCvatD2ynY+fmng0
ddffNCrmoWdXbLG8b0i5OCkCMqvT75ayzVQeQZi+Lv9MrLJMgm/pUKQTQGXaLjBI+OZHBLBXelZF
pw7wMKR2Svq/iqfM+7hszpj3EY3uQOIQikdvFF0D8Hrw1IbPT/ZDgzJd9vJkoZTeoD3dx6TaCUQe
DD5LoeEe6N4oqGEW1YirnOYQNLWj/ogv3uE4OhDFtVD1kXDvt/ZV2ysFVNs6oQIIvhrq8a+L9V1j
rWOWzEuDbX6P+Q+AfX+a88aXgeBmqQLvx5OlidZc/tS2POY0aUL++i3jUwMycfYzLqn4u6Mzz0VH
Kx5FhpYiMOoyiFHr29LuAEv9RBopSQLUVBYyeAbj8RhC92fv4IZFiefy7UO+tIVJIiJpUdap/37g
R7F37bYnz63k+XVdFAEMZ9fkafQ65fgrSomofxWCs8kfyShz9A5n6B2dEYRbvtE/HFujDtJTU3I0
jjE2h+UvhSv8goZffMOUJqdUXnFJOjC0KuA9upY9jNS7wIqcrdaqtMgcW54VBXmylsDOCldOIH/0
fo28ugn2QxLFE4ZcfwWXjHiYp0wXKev1hq1MOeHEmN162SzS8KYRkKiv64D+uW46Uwx0cQkhPUC4
IXTyyxOUJ8btvCOybTPOnyZhy5ft9E1ECL9QhHu3VL7imT5gJBiVwGYXgm8GqQGV6VkUrzLF1KfY
Kn3uKzzTTdtGP2AQFEKnhgZVrnrPth+J++Fn68cFtVzsQcJiOFeYtAxbY3qLX53HcjVBLMzyJq8D
fi+G+DTqEiCRHtJkEPC/Sc15wH65etVrczsIH5FNhWDe1Xfq0jTn6mO+Spz2S/+yxPUtpCin/MJl
ohKGzBQsT++W0VjsJlpRqFGGag8YmRYyYAhzl/w1z1cRopUm/3Itr5l6a+fUzxZscJtYk1eKZXSN
QSJFdqlumwbNHPvm9W5bZ+QwvTWf0TtEbQZZ9x/XDvH5X9HKvz2uaZc9AvgDa7zxM8OCS3ezeLXV
W4gyb62lVMgjsegedymR7vBGCAynrw409U3vPN3PAoahmdXC3wtJmvCmNc0Nke9sbRHX/FXLi/2W
fxxufahb5TT2oY9qBU2heMjooc7Kmm+8m35LV8RDbiaAbMbZqAIv7Mdr42tRf+2irKWc7mGdz2Bd
ESZQ56TWKRKwu+A2DgUmc5L2Tzre+0NOoqZXmXDKXmK05qQup00aisPCRRUH7KpekhVWdRPW9yOi
yTm7QZ5gB5xnEFBJ5UcBKZX3bxokFVo8+YfUS6aV55CYRDzrNSVbYj5M4EYNG4m/BEoC/SUo21DU
yq7W9Cb739MDdJouyUmCp7RQGQbsq8ZGRgkWE2DfXuAGTv63xrpAeV+uf5M7I7y4D4mwArQEfwid
IyTvWUr5rHPFcooadpcV0SwE3WnpHGNeIo1pwKZ0mE1rnH/382ObCzdP/4B/XnGn0AeKQYb+4ZZE
kPFaQhdvkgq5dhBGLseh3NzRyX/D0/b0+dl7UQwlZE2EUWCZ8ALgXezER1wFtDaCm7nor2Og3tJQ
ttjd1yisdk1bpUm/2hc02Io839sk9uT2tbc0FYz8xUKsHak55eT+FzjAD9jMoEWhfX6UXgP1EMdk
QLO8JsHJDpE/cHnBgV54W17oIxvT/KoyesdW1zhxyy4VnZzcRjC7FE2uy3dWAwnws8R112LltpU/
zAq/TGmkjmO/J1RGowIwvWQriGF9WdmYT3mctMS/u70Gljf6zVYgRIbUf7Me7fXmpWibIHiDi3SJ
7EKC62+R1fLG/02Qy72MtxeNxlIx3wAfEi24iE/Qt4PxHmtMRCCyNwsCvt913cjr7NA6hQqHPFnz
toui4+ps1sbL3bjMtSsS8tUcuG2r8gdI5bPBHDqN+ZIXJ73VK68al/oDwlwuFFri9ZsOZVLsMhIF
r3FceR/0xTIsifr9tf8DOKQkeyLJbP5Vn60vrEI+oXsPENLk3WfIh2uwJr/tgl0/RLCr+Q6w3fpZ
O5h0pHpYVDvr5RWlQ6IU7V8sUmAURZfiejbFptOWDYlhyC/GPuR3Rw1RYpuWKplDnzppvFWGuJxW
vZQfBzqTfOng9wdUV135mSvuB3vqAwtmogdJFnd1lhWoMyys9K+6jpuK5T1j/8FgbVUANjLr8rb0
AP5YRH8TAQTo9JuvpQK0NHRWtKX9DAcEThtpz7VDDdMMuRRWHl2IHq8bsSncCxlhF0u1KEZSOODG
vFbyV6YiptNabD81wTeVyZMsLofRYCp454TlTsTbwVnEHIsFJ+pIKBEAzQDVOo5wLUw9ih5M1+p2
4JIGhb3V5N99FXZ4A47DP5ia441rvlHqY8H3EGaXa2m2HNbnqzGgMIm9IHe7lYK7zthFPMKfXu2a
BWsZOsJLLnTk98EPxYFRxaH29dwGwKir4GCO01kGInga6nhaqN94ss7tlO+cZSAt0tdEiOGOg/b3
At36qfLS0ngjiKL9Pj8Vr6gdj6cnDTzXI0xNyDtBLwO/ysv73Vp87Z07VnzkPQkSiaWRKvJjypcL
v19Pbd/NspWWHgdBxCcgeZ87c7Y478j5M7rwV+On2g5Yxjirs2u6MD7bBZCTVTgxnsqRfUGqQq7V
I/osm3wcOAM9RJbpKRCsL7+naI7b9HYf/ewsTsK1p/ffOB40xh0pz/O4E/I3q4tnwg8LT43meC5/
dazfpTvK9OP+fdtnfM7wFRLTmarbT8FlUYUgZzdL9FLobPMM7QsAwshrLUSla1hhU3qaatTWiXEc
j9NSmBL8cpg2j3XnJzsszNN3tqcYHEeco2AebMRpW7bwLvFudvwGX3FPyyNC/7aAAeZ3v0+5xxih
Fc6S8iDNnzs3CswHvTL0ntWsWAryXcWUU5SwvgKDxskH3icYGSKvO0c8JhppeWIux6m6iT8WKNf8
5TZhH6ZSqLz5ksAl7kdKP4elRR5nodg+mwmh6ti8WDhljB93xN2Hjax9SQ/plyxfKrmWqR/ESBWI
hV8NhjpsGweSGDT2x02tFuhgKrOzFJ9Y/9KdZF2VlZSTSTnDReERI4fn++yPT0drUYY70HS2c3Kg
/38b+dM7nPgJPoFt2xkpEKfmBAuCVUUzG9n/WHSwT3yYZMKgbVLzj5/gOvoinDmtjuYkjTPWxVNj
r2BNYODE8lT32SPSSXXDKa2FW1AUW3ulcmVWi31tdZaKq2ex5NsY/Fd811ejDdGvKO65xHZxOdOF
IeWsOC/GE9G80RZDQlV+11GspueiLB4zH7U/lz04EMXuysKHdLTSL/3EQuD6DevS4Tb8lW+UBC3a
uydqSjRztTsF7l8mK+nBZGMNnyCtQ4Z44yJYQ1bF0tBfLeVZ/0ynGFyBvIDpdiWEYE2BVExwUVLY
evV0yrY07gWLoMw7WwG5VlQRhRJB/Rt7U2eefsM0A0gudtBY7ecMgO0Ptx3ZWIhv6DSmnxqtFNtP
oNpIxR/7H+qRJxpiLPMFLM6mTFJD+CF2Fu748Z2oelUQ2kTPJCiGYShOdC9+6dg0jY0kq4m0pZeu
WgCJljlnc2gil28B94bNHKaGGosiBQRGAKgYgwKX7ml+Ty9nr8a8A55eZoN21fQVa1jqGsPTOZur
+dVjunG301D4rPo2cum1pcgJh2u1mxPjx+s90GcZuB2eCfA+O/Zud6HMAbeL/yY7pZqrGYvsChrI
inplEr/CstBe1eQNzO8CF6bItKvcxnoMlrvqhF0MSAkjFx5nrXaha9Q0T+n8NJgnCpl7ougmZVJg
Uic+jr5Zam0ubSYN2ZQfH/G3NGhddnjPRbi+iS1sSjlduRm80XEKqZ78hSf2YVfkjx8W2XIVnJvk
EQRFLjfwV5iGoAFAU82Yvhaw7lquGR/Po82c3pmrGg6coMryoqf5oXCtscaqJeWU+HB9UjBBUjts
QZEa9cT9+X8lOIBVnN/Pl6tavN7Dc4DIeml0arZg6kN86kRYJUuU1qDnung0nJjr7Lkp8VozRn0D
n+Bta5Xtz2y5P829dnPSp88NC/uJ8G4iqxSvj3lTSZDSddbXzsSkYihQSCbYHwOZRfC4ZjPTV6YQ
uLK9sjiTnAPFi8GpL3MCqfQhCk1OITHPs3MOBLO96q6vEQnw37TOiqW1CVkXQ1JFsC6Z2YN8f0fM
bcs10UHcurgVaIJkrzNWfBEFcgZlqd5qnyZcsekk4NT8agcyZO6/toS+cF/dYDI2VGYhvDPae0jz
152VNcPaqb+Tx6hJyQgA8eMUxcqAH09DjRkFTxADn7ds8EKwdU656pCJza9Zm9iItBnhk5DJgARC
a66TckpDC6R+srxVrogD1V1WnZqYVpQok3wosLJCKv0PVGlX5Eg7QHWLwRbRVrOEk8fnXk8d+OLI
hS16pgWOL4PQk5D2Zh1/Eg07+ofX0d/9pIEqob+kH3k3BhdQtV5Pvp2CtZ9pSWXOS/jNg/NcGypp
Zo0CLf6sTQsYGOoWkyJjUB6+9wPODhRLu9Jb57zQ3cggwprK9KdgFKAC04X9eVwvoKOFb7LHtOpO
SHuWJ912SBYTm5yGBdLyHX6X03vIfwv9EGoU+ocgu8gLt0uaw3VfIOG+ctsAvQBDO4ISLQwn89L5
MXZW3upDfE1QyqxmVW87Bf5bvZRvL6JTaFb6sBs+yv+XDsj6FFyDvtBcvT3LD1SxfQ14uW9MnBIe
K68I3WGrr9y2tBT6uFHq2Ksr8Sff9k6CFvxhL2r8yoxsAKwqpKVqybCVJS3Sd5d6JUmj3ndnKtyg
ryqy66mYU194AtejKnO3hwEn3G0MmjdO3Eu9g0hS3gFUZS4E/ZfaNfmw0e1mWZUMDZ93Gqhx1npf
dug51b0BRR0/BbDRUOHB0KK1qoolZ9v2U2+xGSiNFTVdxE+i+ecFYpGXJLm88Nk0fu7YAtNWB3Ql
qk+K3xtGU0FkZExKIFDmzEyk9lzEG1p8N3jyGdhQzUKYQiR0Zi1jhrud+ndPbJaW0ioNZlfdqmSj
pDsieZ7uibE5VlbBvWictUlCfLPPVmIMnaFWiYQgER9by2A17hIRi4AVhUkbxWEWb5y97ysaOWrL
tJnfzXelnKi+URoiDidgVf3U5APsOyPOZ2hYQWJWVg/QPr9eZEh/osm4BmxLthCMyZ4HaAWLFXgb
3vvtCYaolnyW6o2NfkPi+D4sXE6p6BoKzSAAJ6mCozv3sNuSXYxQplwuhetLrJbonZdGkGV5Awqp
ZiFSOk7xenYszzMPeSDNJKBVUcxjuoZb9nj5HEF9pKbhPpy2Xhn+0VGqukE5jP1O8NNRZ1w5Onzr
flSYRksdY065rbbCyoOL4T5D7Jox0EI+j8TIk3hEhObs+H/Kmj/bAqwlxITFTwKg16SeftF4G+wh
H0Wi5VDA2KWccwtsM6uWcG3jxyGVyt6c55ISpsYy6hg6K4b41EJjqsgAmFcwONuOd+nNqr4D6B1Z
5iAOOeeqCn6j+h/kFhwYSyxxbnVL4aXH9fGcYC8fjt7vLqXNgy1paUXqZuMDMFNWDx5aphq218wE
U2Djxf9kEbtWxW33TrbcWRyRO5fdkQuiIUMxG9QpnrmqCM0WXrmunrsZZVkFanrQYu5zFYY/OxbW
5kRFo73/ZbZQqYfy6q7RU4eq7Je9F9V3TkUZmtFwI7nkFiFPoLYfWWOAeAg/FND1CBA7/Ag87yib
HPhX91SLtw0GqrMXv0L68Mn5Mjtz+W5MvrfIGz5RRL/rdqns1B+YOmQe7s6ITGgiWKq+XEUp3+sX
R6AzYy0tjH+st+F1mBnAXtOvMhLPK94bV1nxUKwIvvQvIAE/fMvV4e9NgdmmBZQXgsBkzCYLXxpt
GnNP3FUg3xovcDPdSQzGzmSts0U0Nzht8rhydINnagO14upfhndnVur8fc4g07JPMHcdhTlJdOY8
FQdnl+ggT3ZqfCcwvqqpxat5DiKHGJ4+2r9I/fUMkwfcaQ/CEwaCn57X3jxSd8FYGtPfUHkX3f8X
vChdJV0LvwvfrLa2EZH/jMw8mEyTBLJC9HxyKJY3CLFYHYwTIlwJiREKGRlyRrjvI07YIXf+8Npm
8di9XMrKQDiW6jcyo9QSy1X1oq0RvdJthF47AIcA2y8LATfPJ2P/oCL6VQdl+R4Dqww3J0WeenAk
Pl8uN5COk2qYyuGoUiftOjhWx+SMbi2DT5qBCgBVomsWPhCwAkneZYWgbqmTu5PLbzy1IsKH5JG2
Wn2ZAzYe9j4taiHir+Mt+tSdzWkgQ96Wd19HLLOPAcvAzgHfhZB33wavtSwl8P7B1sf+8EuxQlAN
q7ftdKJSF1WSdRSLDR6O0WHZArebi5cfXQ4MB4XyiJ/qG5SQye4xwMBloD5zTvZdhp0FRJUpm2Ts
ME6OI8zoInpecw4GSEa3NmCYXWlXMdH7Gfx2IK4s/Q1zZIHNO0pzGW0Ik1/hNyqX3btLf9FAsom7
A8B2rOBjpdhLddYiYZc8IsCBlxibDUyoyjxxG1DL/DfBwyVanUw2GYpeTb1kItvvWqt9fcED35yU
o4KOyAPAsQhY2YZxe5JztMWHX1e1mU6UHLNeV94ZOS91yqMsAJU1Qyxz+FGFrtwxQawkgYj9otjS
nJgU86LHqFxrim26MY5KQZzcPQ1sdbfCFBO2RwOYtNHEEeCDYDKTRTZt9aHogvlcWAoufU+oOTmB
dEn0h6haKtFbhfcHOs+iE1FaVZCiKoXkLPIVWO1y/ptJSrymbS5Uvv652UfZgdg/6XWfK7SFFkQM
4D6G610Kk5/0yS3Da2W6Xo2dQ49/h3HOvFaAGxx26Nmbw1o9kazZGFhjq4BeGkiZLqoXQQRykHaf
+auP0UlIlM9QhmYE82b1bfOLFvS6+rJmXpqzNyUvhNa7v4SZ1kHVqlTVmwh6PZ56+2eAj2wOrga0
ClVus0Y2ooOE4YRKfIWFhJdDBmI5kV0v2lMvO2Eergkt2zJKzKZMyP+4lNbu/FeDQnFbR6t/Pmzt
sJfuSZAw2Tua3YqZidqv3U8yiG/zOI5q926vcParRtzcp9yluqcACA53gZ29O+2laxz6+V+2BlVt
3KWKIo8fKZOh1zA2+hyKaXniIKS6o59cRah64Hpp64ejKzHoFL8wQIrmI44wKtM104wz5sDOAUTK
6Nbun0WzSvnKlD33oYNBtrHL7Dy870j8y48cf5KoPe0wcJTnroDkv3e0MLeEO4gEeOi6sRSvJb4R
ehP028cD8GolXhL1TKjmdFSEp2czF1QXaSKxX0QLbnShuIqsgo/6bme2YLw50kVb+Ytm6VAPehpQ
aR4Hjsuzj5ikzfYIZJklkPWmPGh2XotLKAMUw87neH4LY6huL3NFata4r/6wcZSwLwvaMVxf8YZ3
a0yUap3htiWYDrr5eJPHNkTL/J6J97/26VuP0+iXyvdH3gLrAdHJquHIQbdYTNsJB/TC5CUuGgdH
QXjknGXmHetb4sNXnn7buKEitX0/7K+MB+PvebzxpqWFnYmbO8UzYrzwiMQZq/PsOw0TM6BA3MrQ
vwPlt9qC8JVqlj4INAkl+hFtpOhP+mLQ6uh15ZkEkOFxxOkOhuF5CFqz63xuw9gvOybr/i2lwcUH
AplPjZCy5LwIXGnxBPtCeQLzTcHfp62VN8XYqB1yJfIAHSMeSE3Dx4MO/x1kB3KaQQd2XBwl81Ao
S8Ye9LtR9ZCcw/Rq8Slw+TP4Vl3oBXed0+63slkRdGQYxkWCeSFUXHZFVunZVN2HO/jiPS9Zw+o1
irEWLKHmUWy+pGb6Z3XuRyZthl10otWW/6M6HY2qfnMXbUcVGtg4MIxrS5T3cuy2vLPqGthHVCP/
rewmz5hEEP8ABVBblp+JfQekggjIRYoBcDOPlNmkZe15Pah28SvE3VjMEuc4EE78XBslWatO8ACN
TEvT2irRNu+wWCvJ/bYb4lNqjvcuLbV/svGEHmdZh9fwp71wguLGZi76KNOTSZIu4uuF2Id1++Rw
kr63nPFvU+qNUUUPtbO7Dqo7eUhZLXWwdbd3b7LLf12NlOcvK9ya2HzL063NvToKwbajbw80TsTu
b2G6lQJ0hnJSVMxrXUTHcCuTFQcIjLL5VTaMc+yp2oS2ICbVMlEi1S9uzjopKuDhQhtgAq9DlAfx
VuqlDXe9dhKNtBmFsHazEuH9TMsRQ9bWsWIC82tdW1Kp6FwJSIZjzJ+BPC/8g9w+tSXvqmx00Ncj
v975isHAYmFV6qfU2bnSIEQvgzODSxRH/M81fdYJyWq1wY4Vw2JyHVkOkRBNLoLO7PNBLNTp7kgh
0N6HfFQCRHaerq11ZdNFHnv3lQ6KuUmbnrZvDMRF/nagTuWW4m3fjiyG2fSjZhBF6UGhUA5JOzb7
reoUZS+BZ+kDn9oY08FkWqzUykXhVX60vBCFeEVTdAMRaejYwxzg41lTNjXrn99pVDlw8Ko/yeLF
2srawt0flymWHn8qDWBa0brlHW4Ws1Y0XUY20Y8z8a0X+mlFOe2ajRsFBhF3S3QSSiOnjiqg+/uQ
+oIXL1gqjcUoEYHuSZg+rBaI8CVmeFqxtSHMaSoiNPPXA1QL4hc0lb0HKS8T4fWj430FIJc6dOK2
6ivWc1R7GXkkzCanNCCa2NGccBk7+bEVSa8/0V5ZJweaNd05xg0iWsCIfdMkxi57zMIlsIxEbQBo
+VAsBYOLsjNpRv8n7XNzR5qkCsCzKjt91ryI6Dt8JkYqWXg465VtsgKUz61y4qXTSM3iZYtI2Kzs
qXDbHT10ay36dKfxpDb7Lcz3spmTyxJTxBpmmrxmyAB/CFlJirAewCvAvNb9nMe5ayG94Q1aj/uh
LCt4JFKajzTCs0gREyjZDa5noIiyILeunltmSnC2FeNkg0TUtQ5jiwAru/Z4LBNVzgzk0+kQvk3q
ix0343H/jXo/e3ibwRyflD7SabK9U9l5vS/eX1ngX5ukt0C8YhsfLAvNspIzRg1NvpyprPORqkKw
lW+zA0hJDce+D+6uQUXwgqunfR5yI5cPVcifpSG86ByjoagC6h0Ww/SVZqYJyJc8wIPmxwot3v7p
+75bJRHj18oq6uK553j9HafCm/3BZUuTAlXp/NItitjWlfKjcYjn6WfU40wFbVYMwEca282vNf2H
JkmJALaJZfNZiN0EDk+YTRHEcR/Vezi/U8upwG9ulgjPpDCjJo4vpbiUXPCJMUc5hVHFPgVeyPWW
pspjGMY2/ihaUTPQCSrHDFwrHienC9X0xA4kqJIV/j3k1fNeohLkx8k1xCHN+VAFtdFKYnBb+adO
Bt6cIRm2PrMlnBTeO1zFHjrrWg4oHD7xxafGrXPqBCfnyHgyo+fKArQLm0FqF3IbdqPTx2rRFZIf
IyLvo3xfToM2UKdpCRg5ZizNb9+YnGbomqy4LvHssD0NHqrIkOsldjckPHbbr5bnlI06TuSgucwW
0WUvD2vn3pidWMTaBFW9CaaCfQwaDJSeIdujvjzD/2hVAIOKm8v9gTlbUYkbWZKsiKszXxG8m28m
PDYhU69aEGfTlmJBZ6DE5Ok0fEGDJz0kbVelvob8EiC/wdFqplhRXxF+G5bYLmKRlyZweZ2L4037
KQNkAFB/uyd7dzXatjts72ijy+RwlO8C+65BXyKIxXu3eumJTQXbqjrM6YTbLLfntdhDNK94o3EM
q17jwPDZwXRiLTcAqtIRd+C1Va/LdY+XRSUXOjCCnTiECvDnvb2Fxew2r4qgCYAnNlFsMHInjIpo
ljxaLHc4pgPEpoDzJdE2+yw+uNinhXUcZLu7DOyIMeqcwAkxcAzL8iF6EK8gQKEjGiT//EEF1FGY
Sd664A6zoLJOVm7GGeI3j0+POHGZsqf7w9fdYcWP0gzD2h2lsiWpJwhGAR79e3vIHljnMpO7bj95
WGCVhci/9Q5DOEgMpyIIuVa4dOb1IshrBByJoq00fdQKzn1BEnP3OVTu6uZiLYYsacjky06TzCS+
8kijdpDMQxU0yjUEiJxchFIsQNMvsCm7r2Zk6Qj4WHcuAZ7HQ8sMyorFEinX9fuVl/BC54luvO+5
CFJ+YbuwapCuIDkndJygfmn4XsG3/I0SDbDnsHzIaPMmgV2CwCQ5ey3M3wNomkmxH7LyMJlydYfu
PtLDHsB79wR2oTyVI05fMwczXmrLonXt0GG7bPJ+AJto2JkI0ZS5VCuVW7iBsvXnzckAs8tDgaZS
Nm1s0XFZKXrM/xLYybKAm3PX595RMeXDKNUVzaUi3GyIfeltkvaxh5XBA7N3BIzQnwuvswxQDQqB
kVTew0UVefZVYd5bHxePrgzULtLJkMtIPSboOnvSEeIqu6eUfuIuKY1SVMBCaNIhNcwAEZ8DzHWU
Epg3+eK+cnJzYCq3chB95vXYrrNxJ0putQ5YIC7Fexpy3nXKlvHByP1TuQbD6mdzMClq0bE/exGC
7+IsaXhw1DCiEBXInwZX9Im5Mt/Lvy1FYM/G7VFjav5yW2rCEWHaxxrLwUgvX63012yEZl2N663p
n+fx7+V5UXLlKi4CGlaJIuKOlGW8Htob42k8DQl+6kTFvP0pSeG8MZi+mINFKtNtomOC6UpUKrTQ
NdpJqtTkOir5rpmwZ6hPS5q3pQtDEDVcC3TOF7cSNMi0tykBhrjCMKVc6+lWKUV9qRi1WkaxKojR
sQA4EbPLdLpGZvbWY1tey7ZBhp/bLCco7SRJ64wYwpUEce+QIGV+Pg8hLmylR90DhhqsboPcG8re
Ytjo/NfZ1dMwSPrvh5kiu00y8rsjo+EliRnvU4CUCzLWSxbAKkMDXMBnyvWprG6ERe+eN5N8Ekya
cLHvWScCEfhyQtqQ+KvrmFqWLxJ11gd4CbZkmMhRzbj4vHUlmSECiUHca5+43j51EinaIrWBbg0S
jpDcnPQCaZ405D/v/ozE8ZqmYzYs5iHtkw/iTC4OLi2Nq2pN+jNtR8DLDkbJ2OAG7YRz66Kdbecq
IfXEo7nIMIUlXlF6UjeRqWJfm8o/DZ3L/eL3mXtJ3wSEHpGcDLH6LqZ9o4PBpmg9jE2RyMi6ZTKi
xgab70OTpSCDk05FjR6v1174GJNVwOYlPixir4mnwW9SBJI1PxlD41z2S5Z14NOm6PZvJSrzhV0O
Or4IpfXZI9dKuMXzZo3hV8UDLwwt3rcge5HZ1/KWcped2PBXNaJEgb8J/nZrcEz0XQ12x3GpNpf6
H+q5jvxGc6OZg1F0fpwpVGFD2NHXqxUXv07Wgj9o195D8aMou7/0uboifH/Pw4ZWPNr/Svd+1/dk
u50eDBq5hLfOxVxsM8+t/+i8e4G8KpKVe9vFxWoUyTI0IwAKqyNRwqMlyHBrgzeS9JbnYQMUY+8p
N6UPSz4Y8MDEso8cLA4/lg3XTEGZDzq0vCthYFTcpzY9Aevxn/fMVirUK7myReDxFOfEQaolPt2k
eg/iZ7piERXKwaAAitVv2wjDCo10ZXxVzom/zj/fHl/We6pajRg69QD46TPcc8IJl9rDTupy+9JF
P4DrtVHYB4UXd/7Z2Bo1fSTqQpLWNEiDDs8PrISd5OLaanGVm0dHysSIuiok9+OKdZnpB+Lwd6t7
LK0WbEURqSbauT27HwwBaWpPLLR98QxG/i645bioMzXq66kwk+NtO2VMde4sEhNuERT9wnN0eHcd
edo+mpttolQlX4lytFKYs9qCfje46jB3D6PKiNFDv38pNEz5Zj25STWiEs3ZKoZ9XwGPI+dDV6bX
G0lOdw2OgF0060N6QBOia4Gj5pnRN2QLIH99sHIn/LF2U8CvbGzEDONmJ7N8VTk5YiMouabcMMBL
gSu0diycd4Sp6CTC5deAxrnzGCjZ0klfZP0+GPwru5BXk5pOOK55F2D2NP/Q7JWLUHl1G9sZFz3O
JBeww1g20WsvECT2S1fMsX/ah0zundDvddgptkSvu/BXuvf9B5Y3cb5986eTzTA0LXuXxeC8M2vI
BywdeOBedQm/F+TgeeoRtaIeL3LFxNUxghUSi3elHY8W3ESwP1GmsR8T9Ztu0cMc/D2va1bl/xQe
tKewKeqTxdCSuzR8scMaRmIoQFjLx7rhBdNNlppc69LeZwUybraQoy7nkVhCGVGel+aAzpGchbZ2
Lu1Z+/GXAThVwog+LgQGorzdjlC3s2dyuJdCF0ICDdweM1b6AAJBZf7N1ic7QEAtWdh6e5GOdfBM
m5wNRxNfaKNPzmQzb3SBXWWI0SwezXIljorWcKwei+IOWCge3cj1fvDNA6zd7lvfrJiiUtf/ycp2
g7b42wiatW57tIMqVa+/bfoVBFkVgwhPjysAwiVM0r5oGx5ZBlRPf3pr7XC+yxddYUIeUkKRqtz0
oS8C/J8mnba5IzWGmbY+fOJiOVTPsrdc6VyZs+p9lcQVNOtANduIadSjkomrrc121oC+8mIQXDTT
ujavXM+gZBvEqlAxhOoCyd+LCPwafKgjCRqcuXdpPytPy7cVyv80NuA+O4viACA5AaLaJl28kkwW
vM43alyIu0+S//eRZ3MSajeDd4Ptu7B33R2Fpf9uYTo0SEBPyi4QcrsXVzv0/lDdsJ4cQmlvOxsw
o6/wsYXCVRzDASoLjG39QoV739uVbb2uClElro/zCLA6s9GrXvzUbDHe8pxjm8kGFG7XGzFoOM3W
ykO8iuQShh+jo3KamzOtKk0Q4jgvq+qivmw5ld1WbkuwbEju2tMU19kbodoqoCS6FlJ0RyW2gq4m
l8DjsDukMlieM5rOhyaC2Iu+iC7hJG7uCAnrMZRc8USVP1QAbK6UAA5j+/F+eN2PtQLoKVjcCEUp
aQWbiTs5wRfae8NemCNCP9V9yDt2qQxvF5HTnVHkp91NOraKD3YwAJTCSngsB6Th5qSUbLVm+O2/
zDTph/hcYBQWtRBrjXQPl1I3wE9jzqtTnMwM/Itj22RdN+MrYwWFnVLarEFQ5MqpAzm5eaCJE1X9
BhDFrRnQsgT+WC3QXYyZlwX21VWqLECDD4ANjuoZ0foPslQf9lR8yrzEmxdJHQ4qa2HiOyYO/ydh
kKxmLpvFboS2Ygj9qRCpvaHMvjSvuprHb48HDVMprML5+8PPdI48FY+OkT1cArsSdNo9Pwlckskm
zr2+cXv+nOoAK0ayXwY44kw2l4Ih9V8eDnlaZzBXfsdY2/N5J8N/5aNP2qbSrMvJtwt0QR8c6tFZ
migB88hvMGLp5tyCu9xQiJzh0htR1DQY5N42SmXJVzHOE6bc2hTmgmoHyLzMRJ84KblZKlz8ZLf1
LS15TBLfgEawvsQ/zV68nZ9ydEplz3QmVWM38kVGakwKUii6NPOpeo6u8JMvPguCBnrmLh2pjpdh
jPTTB7WZhNVSTVTsGffeCLY3V3iNCuTpAoF7U+4gVNZLbCQ3pyAyZYXhe2pRU/BgxLx+E+xRWFD6
Ekc7WxT32DhK+EZiTNx/vsSlkagmdp+YltLeHSXtLVqofnwLDAdml8/ydra16tKT5B/wqTvWkt+T
2eDYm4ICC1AGQ8OmcsSAQgmzFasV+afauukDSiHjpEzvGT6Z+oRte46tNP0cMOTGc8WxAau99+zJ
V3ZND9YlA03XUQ1JCIwtiIbRc02iZeanN5t8Uz5eHZPJa8yEQhz7BXlS+mYQlYM/Brd5Rw3hniMI
xglfm6B0j+fGHaPHfHJKH90JIqMFNfvzogQt/VLIAifsYKbD06ClvijoGc+x713bpByouvAcSbdO
0TIM41dHIBw1swGCUU0NtJiAuD5H0d0SxW7OM2diKC8vm9+vZ3w1wMFqWsH+dYsvrylyErS+3HO3
h2GaZKswMIcRC/y/MRBg3TuVvyOLzxjSG1xPxuv8B6jGUTmEMuHpkmyapVFMQyrYiEYpWq7yWns8
HZ1OGyrRNWONqg1pXIMQg8lpMHsokOKBn7oFWAdsgknQkM17zYXscjWdhWpijmpdSDMDj9b7ewdl
GdrNhRAT0NaZauPrg5Imkj/Wxl+3cp6Jdl3nLmsb4p601hAtjV6RWnpIF9KQZL/TxR7OdaM/vk+N
EOaz67w5jiFyXPdCq1qCWwFGs9DpvtcxaQQGV4FHgy+0hxrrq1y9+cQylEMG0JUww1bmNF9PfiJh
ZjBB/vu0Wtnh3PbRf+t9RipveJq/swxgRZe7cCxxj5pDD9Hg29pNAktlqUVVsoLTTZf1KorMmmr7
wlXMtVKUthTqX4lqSgxNqnCPgSef5nH+MGSudK5PFUYahK86N1bQobl+bf7XuEWIdHx9mKWDbU1w
Ul2Yf8Atrk7EuaJuoZ+SDgnm6JMJENjRjPU5Y8qoH9MgfAf7Sb4pvrdv7F3h70LZpu/WNeMrDgTo
y9hOy2q5Ku5aeYWN58EtCqwcLJpyDq01x/chIpPN0tJsK3UTyYViqMvatVWSCnXTfGofoipAoN7m
DnRlj5Y=
`protect end_protected
