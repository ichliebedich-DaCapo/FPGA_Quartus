-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yn5ft9S/JT09qrQklG7NEDQ678Wf6qOCeTORAixckBz3hyfJ7CMIiuaChWuQkTwXDpU8kOXV/N9u
TC9NBKd04Jv8QjJuMkfpAk443s0NNCdxKcVRg/7vW4ySRxbJr8LwK1XuC5PkjWVcJKzUtVBY7xGZ
7a2VkEurecYsr3/7PRi8LxNcg3Gsu2s0s295qPQ7DNfJo/cw6lheEqtIbl73hzM+hanyAi0PDfWr
2Gz48so3XhIwXzqQJVht9zHcewNVsKWhLUOLS7U0Ht5ycxfLxaSWi0Hi9H7xzwwKxWgRLBj0d/L1
FbDXMj3GQfKxW7ik62a+rWdBS+p77yo15VDW0g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4384)
`protect data_block
IxgXqB8sg1LQbS51xgylpuW2BxBbJdfYZCNY8krRX8jbzhcNdkcsEwqpVHixkQFulNpioH2jcnwR
b4fcBRgKI3ZYGmxeIaL98BurCafvbrd8FIxrrFT16VIXaqO2z15xq7v8mOMdCFmHuFxZ++FSVBwp
mu6VY5JAB9VCGJBrO628I7U0q4BalKIBzjMPlhCWnHsZ1Jth1t5zXe1sFNHrD9HuSKoOP1d9cKuJ
G8udwCVa5Oagf0fiBch/6XgcjVShK7JjBvxGcUTAFL19tdrnKNE6VMDz5Wja1H0CpXi04KUEmJfR
OlAw2VofIaJWFm5f1x9vWS1FBnd43qMbZEIINrKH/nSinl79fAt9n3s2BAPTDW3fTicQKlP2LYAg
b0XvOaIwb3MMmcmpr2/ZsEw7Okqct6Grfc1QUDsDwyiyTet4m3nmge/BI8HaSBOGSO+B0jHf39T9
QGOwi2PjKpX2WHrIC2gFl3tmslD8tR2RampNBAkmh/jH/K9o/WxYU8Tzf1IXle4LARKsAWOtRJqK
rdLavcKVYXbvS79s8JuJ5y1Q08bvejGKb0EqX8liWNE9ciLAPqIi+Edaum+GiwqvCK6U+C00tzRf
IMNu4jf8349+A/iQuL37LwH1vabhA/ouO+WzWSHrE7x4Wvci9zpmpC8TCU9U35MmDiNSGD/VtPz+
XogWU53d+x8AVMotPI/81AFdtBF5r1Qk93/Vz2yMdZ2H5+xuTGL0IHDo672vap40ciF5gDIKq24i
mg2Q+M0bAsGcTocg3TaMJCd2nGg2LYCVNWtGOTQcYOJ2dLlNFv9Y3bZKMpLd3nmECtGfhuDqK5w+
ZJ2rGrYBiZ8eGRps0zE/9H/4xlEy35JlEJl/GjwMHJiOFJZZNbuoFyjFiu+z10N6YIHWeC0GabY7
X1duaS8dQWNnauU6dRvWTlphKDFmasuDsrALwg//Qp+acomvXTSsbTrGz4mZZBJDJRH/Iw2XdxgU
VyQucJnaab64Ko6pw8hizKUiVa5FqHjCHpp5+gjw0qMsaMpy3T2v5rJLA8NWAQ/QUgQfBBuHxFaa
WebE7dqxQT1Sh0mVzI922z44Ma9TPPvLUlHLYQWqLGh/Yh03HH48yuI0NGgCNXoGjh77JM6Z8nOV
4VUtbgLxmNss1mgdpjZxHyLDTDzCg3oy7IVPfRZYLxYLMP4zo8tiEXoVPnjLlT9m4E/w6K4PipZ6
xX6i9IJKYt72UUlvSrMCH1vk/TLrwUsPXUTDk2qgCkYlDwYDNaJRhWh0bSGxAJSfjmFFnrDoYJQu
tpGeIVtpLBT5NPcsipk5m6WgPrgOfVr81dtzx9Jowxsl7oGMidSXgcjbw9N0QTHsINGVG4MlzjIq
ja5EUJgqAXxOKe/ILF5vuHa8fugsc+G9d1B+718H2yjm1fiAMPaY8YqMSY2qmWhnpo1XKbGf+RWC
4LV4BU0pYNp/3nOQjoe0s3afdLfy7TC4MFRhFP07jEtq9akupjoV8wa123aAD89wB61l1dcbjJOc
ij5Ju+Pt6Fo312OINzODGQl2SqpDXvZ/B5Jh4UqyZixFGKmZmp1HZnhCsHTvgBZAZKw+UVQLIkiv
CsLw/Co2bKUzLLskvVPp8JjT/8JpVUDi8KLrPEggMMFWHjuT4ZVoPNKI6ceRWRIQmLsa5Vg9kgRT
+XdOadugFQrSX7UHXQWJ8RqJjaJqbZleSVJYMaR/9eV7Nz0Dp8hb7/nNMqwRCNZ8VotH5W9eiEvP
bjvUCPzcDpRxAKq1uNXgynvd85nwdxnhUfy34ARi8PqCWH0n0hZoosOm7OmXnyQy0mspVspf1VgR
IIhBCmTbppxUMPLo+gLUGIWLNwtueDiuFW8O+AupMTFBOT9rKXWPTFEMcNpc9YAWbjb/k64NESHD
V79A76VbQ7lvDwUbvkgjJUK5HnB9RILe6L60O9NVy2C8ekXnqJmU538WNPureorqb78wf5g74eLT
UrSK+BbBxYaK/XjgMpglaGz0/Ha/0wRgE5mCl6XZYDAxIwsRaAURUZcii7qmL0RUAu3wzLeadIf1
Ewbmj+mOT+DDafCBzW9hpA0FI3k8HnJs6wiWYjwEsC2lQoV/PDkBnR870Py9205cLGDS5E+RyqDV
8sjJZvN6oV62xURD2hQBjDA4M8TczfpW2OGcoAunrQpio9RVM+0sYAm+Cpe9BuJf26HRFWMD4+W0
9M7oNn6qnL/yN4d09MkmJeuM47oSvPbAxkzWDg+Mv1pT07FfZvIPxeX0vkjkPgHYHWahEIvAtcF2
14mK5pXZij1Nhx634J9hkFkD1EQlVi4lhCLNnmxaGw5w8drC+yMIJZkm1hHlkP+ufs7I1OR/FXep
Wg8V3Lk5PlVAhhzkSwQOsaj9spsGpdith5C0MWkpNdHNhvROwzL2Z2AFiSgdYhqjU+q86IetCD2u
SHqQ5OZGbbac9/IJEtye2gfo5SsT9vEco4PLkGPysuzHQjnfqU05rIiFmQ7MUymRy8F1oacsImop
fuX/kL5dsX2oeESlfYUXbS9QsVO/VHC39nurAztCfXJZlYE18a730fWa6AHI6sMwzvraDLyq6vYH
uvNLti1yzAp1oiF4SD2nZ58MdzOSm9uFzRm2Se8mhwF6vP7JjrFsJ5mSYlwl5UuxFwgmcah4ngl3
agkALa9rOjM6UK6OBWcI1X25KzYaONyjFCmWZ9U0AcKIeJzyPYCRAa+r/7zp6ubSw9EfdMJydf9r
fzYSmUi6kUrCvZHaxryEHBMWaO8JmLZXiW2aHR5d4QWwtzJUt7ZD+FC6rr6PMLc5Bi7wK14kh4sJ
xZCZjrX/R2AdJbhWqI5KUjkPKWvTem6HW8v9SycvR8bbsoB27Ho/e+eGCvF/BLQ3lTzHAjryWvFK
Grn5+5i2aVvY55a4pVPOxSgJlwUhrdcjYTjW3A7DlvgA3ozdePHe5VBP6gk178UToiAyzcMC0j/u
aZMnVaDZJb9UWtL8c7u1NFvbSX2miy+sMa/Dhbn9gHbrSabr5paQRtGQ2E3o/irzkkUz5o89zihc
Hjm8muctLhp/uksIzeEv73DKh5x1tprm9AAfuOZ3ar3UsutSNN/NvD4cuoaJ2DVhUHFUBLd8uwOs
GruUWJ3lzwePH/Mu0vmdfaoUHxkzY6NiiH/TwpmWByvJc6ndL8j5G1qfCaTijJxFb4TfAh5OBnZv
rEQh1JxIC5/DMnxFc92CQWywk/107VhLuifcTBJZ2Z9O8mtCPXUN8G3ZpIA1BKk3R3mqrmjfVi4d
SLnimV3OVizy+CUKA2/lngb8Yp3iu1jzQwm1w//ul0utez0wCUcu+WZRwTxzgn7ErptGMOb3OGZI
4k7LY6hrzJD81FtSes8DtTsf9KEX6ubVX9cS6qJyDDYBd8OC2ZYWbIJFM54hwV3KkYiTiqSssGen
3P2ojGlJjEW8U2/tfKA6HNHM2ujvRf8gec/8H+JY1k81WlwrGthn3DVy75hAyCkB+lZq6K/Oc0s1
ey6cewswIwaW3lcQ6ZfNyhqovNy406Uz368Mvw3lJadtouIkNl05Fq8X3nsXunAOF0655wsWAwrj
Mo6z/s5gngwpTUZlB/5pJbiGg0/Ck0/qsuPMFxAJbN1lYSjMr5q4Xrhe4KeLoRZ0HxyCNozZeBbQ
2W7uui01/TuO9ON9YZR3jHG91XNzE2kqysJ+TCU7Kljf6+Xuqn1TcWLQWnI3HoCIm4bkTgPYxBnQ
xA2yWUzPSHX0ZyKurVmBRSGe481lu38FPTA5iVm/nBzxP0YX59O8WBsSSEugYzASV3zWJGPuhWU0
+DP4BqWhpUvmyR3ENqzTblhkHlZumm+S1SkAfXXW5FXswWaVP5+MdY7Jjn/mf+nIOo/Nf8QvIo4R
ZZUJJYOqSfSj1OINSDIMPEKboyn5aazsEHbV2VhLKpLGPXwuKxXDU/dmAJsiOaBDILbCv9LQwt1f
uH0NUnsFtzosudCZxSVGEJPdhJ0yqY/hoDqoP54kePb4salZHpueBpsz0rlTQ4VTsWoqya7aPs+j
pKkbeJ1j8z2h+U3nQ5GNXfKqvuWFAxsDLCaJgibYXEQQZXV8mzgQtgJxmtZabIKgormZaw6Ux+sP
uSHZt9UkvdeQxWwUAlx51QAJ6+eRwOZijPU8ruOEu5M5lWp0sb+4vQYjmIm8RGzehD/zz/W8KwCJ
B70zRnnnkR2cJ39IpklY5BLC1Sb6J8PpZ7RbpwvK9/UGYKYE9vnDu2yru5lLZvtabWdibSZivDm+
A/Ucx0DLBtxai2WSzzKWtFrcj9SGB5vYz46cPfg+9hCNWL+RYMaLI25FL1o2eTslQtRormZ2lgHK
iuDGcteQOpAC42UkCYeny7WAOKOAiMd602PC0R44jHm9z6gQ9r4LNt4UO6Jo0Tt1n+3guZn4FsGo
wETWRHAcmu37I1MJF17lSnzEskl0Qxd3cvw0j2ZkYoJ8uTan0Oyw7eoayu43TL752bQSdLpGhELz
3N5i3VqLB8uOPO2CIL9VbXrCOOGQYwu9dQKk5wPdweDcv3EBzobOT7G9g0I0FEth2CCuWgMjmj6Q
YGtb1HnT0Qwwt9GL7EouYZg2oHgGbMYzvWxG4L9Kh4Q0x5txYDqLhv5WBvvTGT3d3me0xtCk3UTh
JBA/4vysI+MOm3n3bA5ele9pb3ZUDV/RpLV7feiTv30ZJh3V5LP7U/bAWBV/74l+EFheGxIrV57K
NI/qCkz1lj9v47BiPlWv+pmYelkqJoT/hBlEbk5w/B9Mg2WXP+Qbl+9k0toPZZNW/cMElB01SeNy
jWBSWPqUokPV4HHcjZ6tpQfMf+d8HNL8sXgOLE4kO999/0vaSpuUOWcygMK9bQtJcQ55Ya/3vpOX
V4M6R3OKnqn6kFsy+oHgeuJzfbYfehG12ZF/njLkhfXVO/LCcNRXoTsOVfAZJ7nfh9WMAbdv78as
zq6uFFpsq+DQlpMN0T5+DLTs/LujWD2T+NQ0Fb9Cqbzy4I79XCBVywIRWAcL8t5y1PUirpPIP/lI
Cc5insaAWSdLaFp50QtrxgqBAgkcGMl+8IVGBSvHer3yAvms4Wv/4CkvJ9JqFpQxAyTkjGkOSkIK
IDbF/1Uu1fz3487nW0p8o2VDpoWwebPUwEQGQUDPPKBOztChzLhxpjQhty8x28eFd70UzcRyx1x2
uK4mZ/Fg3FuJ84iAfEgyAidn3rt/HBcv21Ne+GZsQOxG//DDjOqXZG/XnO3adBGg1gY0q/AUnpWN
Pw5kX10oUs8KixiTrlDb1KjomTfZNlhhYWQL5HbyXZ6N5pYI5gCkUtmetHFLeTucFesgiIn0nOd2
WgDwG4+RcFU4Qr1e9RNkJ0ko2lkrATdpImElwSA5jN8ZgK+y5oD3IRMaBUY9X1gO8237uxPLEGhX
RfJ5kB0EIWm26VI9E2mAGqkUzmwocBqHqyw+Mqj/0N1ap4qBc4iqjFx4E6RKL20vGC3t0Q5zIOX4
wWWg9gVaEPXj+SHpgJgihXAUVb7HsVVJUwYqsu68eyI80UPlT5d3xCOvbSEKcWU9f3J/jJJZomR4
lj4/0z9Mj7MKsrRKTstg9p8AnUj6qSpxTbH6WcNzNJN18mUKj0UeZp1DiGT4aizYWZycyNniGclQ
Kq5fRgCTj0d/8ZQct8Yl4UvPnaljRXUmrPkAPUMdSm6W7PP1z6HxznA1bDfH8QwEJLW+O7+IH07a
idOme7AOm626RDhPWnSgnZwEcTVWubNsN8QGFTiDYSAfQh8QICqfaNquaj5Jh3XVduPvQ3uh1Zca
jzjsxCxl3Nx3rq31UwZe3YEx27dwDgHb501jidAG6iK+GpnNMq0jNDEnZ/t3lgzD5qM8xA==
`protect end_protected
