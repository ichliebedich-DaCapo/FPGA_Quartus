-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M2ikSe+uODMRsA5+otiA9O0g0g3k532Oh+sx0XNB4OfaE/lPx2GcaYAdrJRNeVtnrmZfXvacsdfC
MydcptXDoGlmMFRSH/ykMsxICvfDfmBX7ulhBlGVc/vp3PxhmYT17qQrYXOiWljEoGr59TN9rErL
a5zn/4H5uCX1H3rFptoxzLxD5PuXjXLxjrji0F9lfhFmQ5+XOkndELtulW89bWFRuPqs0Mx6ztsV
DFinPTHlOsJNkdEmXpM7PddxSSbqwbfFw93mal3EAVug8gI/YuXUAqU0H6smlrfi8eF+rYukaiHK
Ez4ruFA19T7hw2qJOZv4pntPx/vh4GJfHIRXmw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
zmBo/Sv8RnMA6L2A45VEjm1ZushQqwSF0UePR2nk5sVM2ajZ3O8IQ54oAyeGL9+JUICgdChaG6Nk
9Ex3YMN6LgyqTLxdcEjDQqy05hpOL169UPMdDl3urmcCgJj7/C6q5rBaO6Z4vnhwkm4zNgNXrhbj
uXjdeSh26wenQ8svdmJb0k4Sp+88Gl4noa7uvcJ50rfzFYYk7IMe8rBkO6+rc/xi8WyTv9jMXDKS
gOP/0WokzGzumw4XnHj779Pzl9tkOB/p55Rkh9bhgdTxVv0SrM7o1vvtyurdo8jiUv5fhX2SmksY
Dy0LcKRz9//OO8VqJjBilWAlVaUiVTDbqLmIIzNuA5Mf3cDS+3pymnK7LgXx3V4yoeto9Y9gPReH
e0iKqENGaOJarXVCaovHVFpQ10bgm2INXIrgzlokoXAONrOnRea2QooRI0u1h83/aLWCp68BtM+O
JCRaCLAYbLbm/oMSt3OMHp+w8H6GlXdtoPzltQLj4UJ8Lm+pN5l4oh4eSomWq4XmABEwm1XcZP9r
HWuOqobEYR0zETeJ0dSKy7QlhyLjUi3vk3wGzIOMkUF14TtlK5uR0ZBAKpUe0etR7EUPYZ8rlwl/
cZ/ngNVaII2waEb+3JCXNVCLGczD+PR8mJzv/tH4a5DCSnlqhvJnJF7D3bu2rX511c3Mm2kS2cHK
5vOBENozL1XK+7CaJ6S8mx8BqBYU/OppuZ3bx0SLTYcQMTmSgEqxxQLhFDxzJGtHLk/WIA30X2Gj
OhjbXcqHy9WEFqhj/oF19WWRMTFzUwWNPrHAqb339rquy5CzFEgelN/csY+Fv5De9W0urj0DamfY
ShkXp8CbekqPXXmKMzvKfBzejQ+0Q7aS8+f1vXh6+pRG3fuDI8tI9M0EDsixgVU+MXYZxN63I7lg
ESdcBSne+Qi+/v3LcsWl7dYKvX0QH06SfQvxl0IRbtriihzhe28WFwRg6RTxcoEM2H5DPMUbJtFs
5n8V3g0xe+LlSHQT5gsTYJNIQwstVbks6CxsrU6vdlFhTGlPvTLs/zx/9pzUKLn+OrvVD5ZRMwbp
rQ3QhPCJ812fb7ioLwmg319tgK6F5OqYeWgNyEL+W6MUH/OK4bJa8Tq0WKRwB96YqFugr4DGp4H1
kXx8lSR4BIty0tAr3BbBfdfCpDt6YYpxw/yd77VAaPXWxSgT1sV96TxTeaL/6CkCxxtfOgadtM+y
InKqBOcEm3NwOLE7npB1mGWGjaLBuHVr1zGmuIf15uVbo4c4ObpyoyScUFKB4em38SSGFxD6hVeg
bPOyPJ+o4xpflv1Jx+UfFOOFWee3RtRIKjuXn2oqVgXSRnVU7ZQaNSkRSTTGJ0nbLpJw2Q62vI/X
mLeHceHXToGgxo8uuGzHPbIQp38sJWZ9NZDPF1b5qG0U8R14C5khA6apCXgsNHjlqeWnjTe7E+gt
Z+QLGcqbOUHc7JF/hslpdzluKmx4HEwlETJWMZx3Q5wIkaIeXJ8VxTnfWCI+pcxA0kPsgpXv35Kd
mEZjfIkB/y8Z4fBPAbTBQvKxW6OywYn2fmgkA07TO/CSUpAP3qEEdwS6z2aEmyl3XiqrjHtVL34r
bNgINBh4RFoduoEteURU0bGhTfrQ9Z7RPtDq+ElmegDu9iTvhJ9mRrVq0kYuoRRUStI50bTHlK5U
0Jv1WRp23gTKBkRVFSew9P49WMp/TDJ/uXqzCtMA+6cKs97T9bV11nqxz37ViyNnWuO0n2ASKUJ4
5OLhgPjRJy6XENsAEzX/oAM8BVvrgdnYKET/OzoNtHj6yCr5v1gpVUDH9w281jvmZeLy7E47T8bc
8px4bWOylIA46GJlpumyVd9a5bFstmxT2jePGABuHchiRAf/mpxKkMcV8WVDcYfDtJDBmOyHW5Go
hy8ZtcXbxEqbV/Gn9vdaC5DPpLPoWra1J6TJdEJHk9kisTjEHMXqF67FL9yGLqd3G1r+Ga4gpwlU
RXDikwFbzSrLtipVFmAtnatAKtbtgGOvf4KUlk0uUWd1tLjhEvvvrhtb6IqDC20H0iZ3MFUtQLau
FHPd0ySUPNfuu24x22+aT+j93e+CZICOWJaaYxqIwC3D5gydBKvOrB6tmm8j2L9QdeHJs5/rK3dw
4y1NqoB6LqqXNFoSfWvU+LLIo8iYRoy7ecHwB2dx47S4F+1wJBuxcz0RVFMP6zYe5IlOK5r3IL1h
FCSALWdki9poMSHpXTwvruqqV4GEBZPsXAEFzqrVT0plg0Aw96s9K12CJEpSwniAoZU+X/5er328
kKscFiKdajltbhW840uCi45HImK4WKrGmwiI4yeA7skpUa0nx1uufiI5b8jvgc9q60BI+okne066
BfgfXBi1nT5OKgKeHVOVAqjpgSir7ACmBcu1V7sjccOEoTF+tu9Bs73P98c6rIlVWxfpGb04uasO
UdLDyERjtxtGDkpL3IaXAhVYvy/08T9lzdG9cTdFBJ8yJfUJKkzzsD86LD1tbh3J9nFFWL3YAaoQ
PmZihKppshrq5B799kWc7w06Bd/TQrCY0TtXrVjDIibhPwvAjroqtg6TfJG7nr/ZnKo4Dlo7y9gG
/d05FTkzt0hit6GitnS6s30Cfty0tEGcqszG1JTLgfa0Gh9DIM8nDCq5wmD1s6MS+tpcjCOMMGNb
2cHz2wCN2swnKDsP9h26jm58LEWAG4ni0uWpesntorrLUdgFVdnvND9n3P90/QyD/9gp6THVcQsm
7/AhOHFCgPhvtFOFvEPDwdEzKOJcWyT7c7IVZpm7s1mpv/iK9BbJEf8s9SU71wG3hRyaSU6Mk0CP
qEuInmXi6y93zpCPvF61u1sOm3By04ol2bF1k/i+lDVWOK4GTV9jBb/riEwWxKq1b2cm7SIy5Zk9
diKIIFbaG7F7GtzJL8n2nzoz34DasOTKNQFPuxuefU22B1JzG5Gt5wcd2z/LzTSWePHTxDtPQWxy
+onIuPlpc4IOOHFo83u/IFL5sAkpFhjOmz7gPqejqMJQXkq9OXTDcIZOnKZnsL+AKApLHhfYpJmA
vl2O23myHyAhgU8babjQ7XcomEPl3aIATcFb84A2yK2fBM3vlDIM8P6piMgwWkAgX1n+/P081IIP
P1IEBsT8/39FTCxYB2/5OJxC51vTA0fX0R1pdQXY8y7GhuPk47x7icdGOPbHI4HAHp88LY0PtqZ8
VmNSysqAJ+53dxIBCRBG5TWuiD2taLHjPWb2zOinOr0Wc49dcr+fC5enbUmVbSwm0dt7I4olnA/x
aCHbR2cwDamL0IuMiJtvyjyGuyeyH+yoKFz2CUeBAZjGz7GFKubgj4shGiCzQvSCSaJ4SjQB+aQv
0KmXhT4+XCDfyFm9aBetyI24hVPS5k2X/58fFnctXl1oZOfyMAe0dFlNZvt0ZznpCo1jC/5KzZwH
2OIIYlDubQF5dOtMEtfGAVf61cwJSqgEuG2afx3114n1sRsAqkH/C3W2V04D0AgsOnpTDfp53hOt
OMEzef+CRT1UJOhZGl3C4oCmN8gSqCSZmKFGlOgLCaLe3egOknkMTGM/EBS7SHkUSiU55nDjY9zT
FwbgyAjx96Z5pcdWXg5sjKR6yiELeCATXYU2PqzY84mUM0IY54Dl7bFv3EcQ6hTvkjmdr85qp5fr
zaZm+W/4Po4o30LblXO4e58LQa/HF05l59rQifIoSftiLK3NzY1lvkhUqusQ9C1Lm2Lx1VFMK210
NHqij1RnwmO55iKWDw5O1QbJk+bQsY3qkMS97PokXEzVgqyNCmgB3qO5LOwzFAAp2+JqyuNoQlJd
X3lSVXeUpnPVjgbUZNuXL7v6bAQdT6O9wtSRu2wbqCG8eIXOSh2E2AeZv6jHC7jDd/mDAX/QAeKW
Sco6uNuPwDJ8B9I0fANB/mS3yHak/cNwsZ8YoB2SVNYHznZ50pjFRcL08AXnLuC48Cdet+UNDI3R
5cdABQJ1drAoPGM38Qps1ej2XX0Qfxy9Hx3f74eCR1SkeiVKOgC1KpfUGUW8aG/e8FoLf9vLr61f
l9wJLuWl1i9VYYrBsBSAx7jnVgKOOalNKdurvcYTeygSfYh49E+2v9+k2CHU4kvajb1ObpUZNrWE
cojQyHU8d+14TO/ebatjHaQ4z8yK8vEKaT8iDg/XwvVKIMV/Hudviq5MvpxzQcjdOxDOIWYq+D2X
54fygnqcbTvjCKAFoKJo/kXEk9lZ2bZtaB1oiFQyp8BA3MjMeKIhOWuk5q6Kt/hjn9MFUzj8iIE/
lwec2EdMiwJMkcYZnJql1YiPHwvdASjPIFZCGmBlooCRkCGgq5ZEzM/j4eCCRl4baGIV/DwRqAKG
ZezosZkurd8lsGzg84gseQmLmQz3zOxgIrJvrSnAh00u1A1ju5I9Y9UhwQ6V3u0kx0QJ1yoioiWi
ZDQMvL7/4EwNTm0hnYGAd5W2BgoWzbQIC2H4cJQmZddq24J1o+v2dfPrzUUOSkhtm5hPQX1bIDg6
MDPU4mS8ptHMOT4u7YWCyfELzIdt32xFTg0x14LDp5vNoCIfT4aSg2ZtnNcRCLTYU1d7cjJJ+apJ
pxlMms65ZTISNPbs9ed56z8H8Klxm0aqhoQbe9eL+ZDWfNez26114ueixjEjAKZ89Z2mTB8TXbil
5ww2CbWZtO8FgMapfRPGq8mHoS9BBI2sxe2PlED/G/d/o+/namxIKYb0HYScF2nHqqkHKVwAu+GY
AR9oHP1ldQvxlwFu/o6dsJyq6n/tSrqDRi/8zdik/XvEDk09huniwapYhQD5BTsUVUR29HtqFZV/
SBn8cJgfuvU/LWUwR0F+JlvRILFjWdR6XhHx9N1PmU7rEdveGl7mbZ9L31PgtW2Nzy3gpm9EtXND
wsqBUGbM9hsx3M0Oy4NryX232jOjR8MVgsTpoIUL1WIFrF/bzpJB8zRSpKWxxMg2JrIc9JwUKTVZ
oy1ksmnSOaoHCHTaUVexNUp9MUyUrSTFkzGRIYf2nVLtdkzTy2Rqo6H5ERyz/Yp0ovDcUMdMKJmN
vv+k9Cq9ag5mnpUVeVFgoDKpnAln7UyCxBI5nQnnDIxpztnuZfh1aKVCN8Li2ikIKXWRa4nBaqDX
RjywvhmDbk5py2G72Wp97I5qdQmTGaGDEEQ7MB4kEY5DP1tfR0cDki8VsYcnv2G0nhYAXw++D0YY
EJSXniFJQqZQr3sKbJjfUQRb5jVxcQUWgQaQja60N2sK7MiRBg+FTd/awsAu+iN6bygP6LHByQ8J
cG6cFJtGd/ikPK8gzqFmpHA4vBeDKXmw1TaeYRjoPqu8T/SGchiP3VGN6KpKRbnhmIlcOGF40v3j
KCAH796QsMgLLyeyT/zIEpViZCoElqeUAKIAVO1XrpBKNy4MQxMq30vFua6PNjtkAI/K882n9h30
2Vu94WPMDFpNzTSmOu57MOIGVf75q6lGsUUvgk4zQjei6eUr9nCgfVepNvm36b/JhU89u5TkiSxG
i4lnkJ/UMQH4JJNEJM9J3UJhgX4xVbhaBLhYdt/HFASTWYm9fLCVJScad/BH7cTxIl+vtC8WE/mX
vRUkk1E4cKoxmM9iCocQ/jHoIB18xignNH/LTHypoMv6dhZGahIpovDSCvaWIQZ8kcQ4uqPEP5MF
DsioiG3s0/H/GUbbymObJcMBYeTd3EVhKEI0daR4h20/Uwrrxd8NCIWr8RL3VmP6ClNO5Jmd3vpR
nuVuVZ1qthqmPNAburEYuoF2CSrYp+VSNkehHWU/NB84QZnco8CNLN668qRrTVIrEuTXJ7Ll83dx
UNuFvL5uxbYRwGoVMUNj03FxnKD5vi6bYh2D5hPfpuRSmsnCOwfSWRrNfiWQrlAI3IfZUK40ysKC
AkBPHDzTIalyNU7LwDVjJT3mlBubTwy7Qqzcy/Jb3DtIm3/syVmGbAYqtftB7S7eRYuz/+Gn9VCn
hNxxhZ9J1H3JaO6nt3loTVaXHk/1rGMeKZjEzA6zXk8apTFZ6ggs3/5EWAa7Mhxrxvb6cq2sTRMq
cExiud3L1RIxAnFRoevkiTBQHA/iC3c3lMU3sW2s2tEvPfKRtTpSlQNSbFUCSvHEyFzYv/3GdgBS
Kb/pBOJE4xtTmOBwCBmn66XejMFLPGqCKcKc5e3LyhCy8FL4kUt3MGGmyi/rt3faj6BSU5Gav7OM
i0Rc3g0Y8krMGQMAKippPShGtayISy0ChAKurrShoVHIuEaIDryfIR38PoNoCramYRsZOM9lj4+s
FcSgzbiA9UrGbxs6l6i5460VNgkKYaKWWOUZEIgFNQhq3kXxUXFSyLjYXt0JDqI/aLZvZHljUeKo
6ysj+gTgsbMwyNojJmwzjYm4Eehz/ZDA5yECViTaVbHW5NvqP3+BQy9LAn9YP33DGX0sQNHbQ6QB
dIRXQhyXyhiE2nmHnLZJv/yIgfn90tU6Vf2uWJ6TQYfL3isBCHYEPylH3DJBJ3op851dS7U7bFSM
eMsA3uLcrIyKL39F7nopCgFr9KNy2eBbxoaLv/BdEGhi604yrootoWz/g3FOPK7cl/4A43jnHfrA
utwJCntnoZ+5m2rNS8Lr4Nf0M/eCSgagnuLEf+Jg7inP3X763HSysDvsvdjZnVjrafdKnMjY1bso
8s6a+EyYI3FAwCdeSymfesE6XoTFZHJSKlf005EBFq17y7PfC6QvfgwPYXiAzrPn/+2FZ1cAcPqk
W2FvxPnARicRmQXOem3eFHnIxPwJ7gaeEZgaTkBxc5DQvxCquGqHgkuv09hUf0PZtOyTBKoa8Pw+
4XKiInxSfZKO4MesfRzgI7OX2b035FHWK/zVb1kpUNubX9agRmtlLAEJLaV/ZsvMAd64IL3fid3D
TuZlM02g8b9lAwg6LipjUhWJyunrNweCcT81Ai8uBVl52fCfTkwcOPIvLw+5XIdrChcWjinXgAQk
Y+uwVlVzafUs1dDb9O55M3tncZcQJl9yBtfxTDPGGDlqTZspHelAYVeG1QzwM+A6lAlyDrCjm03w
m4mB9tYtwW2lR9ba5LmUed1vi8tI8cfKXAGgOmUIFMp0WPt7rCnKjXGYhQnManNe2XS2ew==
`protect end_protected
