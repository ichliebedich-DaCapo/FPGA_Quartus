-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
j4IKd+x7gqELHWU0HlCEe5LHSFQrQPe2N2Fw1kGGJe9JFiDRIMsomotR/VKCp3T02qTJMPP4FdYo
m5DiFvWqrn9yXGPdOuNQXxT9LhaH4GfbFq1Q7mLIg2P1tsCrJipfpfoNunTxZo6tHEg43Ycib4Fd
bmpTYay5GBCLAFs6dNMThx5wcjcqO6H3VQmKS0y+7zQwgWCZj5IAjcfO1daDP2aYOp5bxQlSMEy7
c3ey1mFz18dMcIxLE+IpH3/46tI/ySz1Xro9hygfbJ+MUxmFoh+lbDtzEExEO91t/BqrTs4rlP8E
0PifgjyCsm+ctshJS7XR661kyUCEX8i1cMsbnA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30800)
`protect data_block
eLUPUIRa20ImW5TxBN+hR6OSR0wEnEF0Pt7thf9gP8gaJlPCOjGBox7e0JPmyB7+2HG6pw/mKS2i
ckiRzkBi2Cy1R/MwBK5bWMjCc53spS06KcRP/w5Jz6mqqLj6afXzS9jkUbmNS2+ATWk2+gLJqByQ
Nuc3GICEYjhDmNi2DxoAkjZTz9XHrJvcjot48RosX/peqacN52YvqAVgeSrh7eGSODcrzP8y2dr1
++Rkp6MhKSzI+wifamlwZ2ydZ9NwQ5NabxHgb0vBRP4yhv6xepFqYLo+sOo/qtLwTDxnJokqdmh2
3bQNvz29BgL0ufLUKZIpDKZi0G+4+ty2sNRwEIjBGTcs89Ckc8grR/6DY6l0PU6YYBSX9tZSQLJa
vK/5SfmbRhpRERDiPx6bkrzrZI4Z5+bWTjEk9sRWd4CtVk2tD1NiCOQ41LGl4qqK9S/NrxSk+g68
5QE2AiWAIqOEYmiOmYDTwtQborkV4SM0pXykvjsitImDaa5CcnvLtAXgCwD6NUkiZQKBNoWRPD1r
uriId4lu8g7wgBtg9W2SlIcQFN9vszH+go55SaSmLhU12l1x4GhVCpb+Ii/kIaK7LjNcihMbWfrN
SiRyCNA8hw2A3+PW9OYK0NdHW+MLhgChqLXhK3Q2gcuEqvCaZtGJ20Aj7R56IMgIknKyuyeTfzMW
DZwvKSRMyMOyyPvnmuNDajXROH/wHiaU4mjjEEo78ohc7OCah17qfB56QL7Y3ypPtq66MPSiVbjV
0SOjMC6kDlllUbj8qceqEyDbW5wmsGPPGtjf0OleGF9gRujDph4nn1MXp1C629KDybHdrvzhtvip
GBmD/agB7vzllFRl8DwVN4k8cHoCUGPK/kISW111Y/F3k7GrhaPjqKIJFiZMOsBcfsozi+4Y34vk
xVZuU9apxMS7mvN2QuEkxmUecVU2sTCBkPkBEffoIARmVi5cC4o2rlhNh1E+29/LSRiy1OkVBRO5
EIkIsJFnkSjNk1C2BqmV6cQol6fkd2h6P3KqyL27dHPILhCeo+T/30gyDL8qh2YfZxvUiZmR+1wI
2HhiRoUAYS1F57UKJ8r4FYKkI6m3i0UbGPXkJnr0wovWztFC816efOPMdaK+lv9uGh2H8x7o49uD
NM6tK7Pl1mV1wlZXgK1kFhqwyHZ9Eo/P2sVW4kfxWEx1zw8wz7Dza3u/oeSqlihIOJ8B/esuipFi
179NXum1enuAzLQv1m+oR1a3PJRrPKIW33xatsq5fJItybg4ClHIE74N3dZD4YhwbYYvV8vv8UuC
uUR+HZheFhbRjV7nvLelvFajaOnqwgQGIIIgD0ZAWo3SlaxjxG1ou09kQ4vT2GLF60Zg6Ji/BSQB
phHlMA67OvCYUA2zT0HLzCXH8hPblRCtxPw2rlNkyYOvQ8odvdl+S/esoWjVKyTeC6BE5Ndp7smO
yxZklGoo64+PqRFlEtA1YTOaw1PwCRZFiNSfmQNbY+PkKhBDM8ZCeYMS3OF1SEqeHasytURSk5ZP
uFJ53c/98cISJM3NOSjgm44QvVRAe2kENysbyPTHZxc/cSjPLhDmg53KE5oBSUY/fniv8Szp1mXi
YzlXX62p2VjayFcJtx3UtWEPLPSgwVPZYu7mBwlpHEKJYbWfJds4DIvDch/OviJ8Z09qKetDTF5z
7CgTAdADiOBlqNq/4JDOGbHS5KS5auNIH2PIb2ihuZe/lLXKbHe7RV/CwaaVxbDGOyam+IM+/smy
711OyclrstmJSe61fUNEc1oDHYXgrLlrUhNUd83M7npqPgV3GvfI45b7GQMxl33Zuaae+EzdtICN
Q5XLSQvEaCah9fxoDQZT2YpaikurN5fcguASc9ULyyFwduVrZPRiYP97f0BAGKjuZnl42ufintoV
hr0sf1AN0v40v4/QnIavdjy15mIcH79itFCzcRZLO+BmiT3m/5dHC/Ep2tauHLcTXExoPiZfIuEG
FmO1lNxlJUKmzT01IFu4uYq2V5yf8wAw3poArap56K8jiFJ2R4D13LgkCD7xHFgn6juqwEi7/oGh
GLoOH9QxTkoBxAqgkCUxeTeEf2bwqeEkMUBE6gauK7eHeWxZuks6S3vVU5M/aDwstMXS7zmnAewB
Pn0V+Qu1/hM9/TMLvfjzjZSeLM4XJQnOS34rHio0wqWNGUiTVwI1xw3iaq8k3BJED1k6kYyCUyDq
QrNvv9VeOI/gD3aA+TckMapjlgxTVVfcsT+wROAg5c7xM9tkZeJulu6dsesKUSq7vqyESshzxj11
HKyKafypmMpTrKunACpv6mWeBMZ3FVZE/j60/TQpS5/3XaDaWFjaAvTskD8FjP8fytdhu7fOXEXO
fw+PePc6DKU+vTLT5vcDoJTKFAdQv2EAq1WEuBbpu68t9GcggFNhB04V+ZgPZv556Pf8ytWlOUfy
9fowWBLkMhQZ66bqZaYbK7jmt09UEdvSLjN1koTJrnAg73PS3aJciEByiyb4JETLsJbqcalPAyrt
jDgmr1LiqPRdIcntuXgLSMhy0qomHsdZsk4rJSRRAsfJyOhRpB5ow/IFNkNUX0wGNjGKOTZ18SOM
+qDH/L62VCkO93OjEu2E5RKoGlnJhwgR2Y7VHyJSWkDwxpPVGbXOxnzR1ObxkPVeYDlGHJ2Sd+uB
1L9QTaQZf/7GO0fZlrqEcBhKmqrAj/tNQSW616YTwsddtbpPuiGEkAk1zGU7TfA3Xq70AHfL8OOx
jEDXD+/r5ylVuyD1wonG/BpBKdX0ItuEQCZhVTsY2U8x8xjqjERIEj6TdJOkug7gAuSdKys1pO6n
svAXdzV3V3kYhBuG7cAUSFhimNKYJk17ns99g0h7U7Ks6vK5sBJtrsg3wD0vXkeNc/sw+0kWPvvZ
I1HH3cKv35QVU4rTXVn7LibvCARnojjIL+aV/Eg3XhpK+JHWo6f66elDaldT2YrDbj+QPO9eTY9Y
sgp8HthpNRx9OK6uSE1kUailngxVjlhwG6GG1MDyZ8XbMJAWL+whA9UcP0m5PoiE8GIyEbcDadEm
4SZwgq15DY7YZsOsq2SJc3hR7iv4AZLPHPPSpUx9rarKZs/hKJDjRunoAcKjMf/eOJiKi+fa1oiZ
fTzKQumH/bv56RZuwPtVRbEsi+n1e8uQjyME/AcT64dWT9eb3/GYQkfgCdzW7+UmIsQhyZJ5MIor
cQn5BnxFRExAchxNQm7W6OHNQasVkdah4qWj6RtDT8rHY4ve6Z69QWhQK4LJLaRSXmfeaQXSAdDm
IzAlhXQ5asmGBZObS8gmV/RinBBTgXF2Nh64o2AVk3ClHeuq8Vd0NTbl7y0zMxBxdxTuyEWriUvC
PPJPAYYS/GQ1SkUirGEdPWDOBfFVA66bwPP5zxZthpWgdMFJRYC0JKC/z55i7TWvdjPhoy6xEyGq
BtdojnSwNpNChA+8D67ezjXBTSxM+QmgpkwL61TEto8peRhAMXJdNCeWTcwv44URy+XrIKtctPUE
OUbfLtetCG6xV2LnnTcJsAK7dJ4V00KHZpXrusxyvPbSnae+mdAriKi86jnMCSlGB2P9OX9n4HNP
kZTvAUs7r4jLo0QhzI0LPj2+yKPomk8YHPi11nevG63W0AewDYCUyzyM/qk3BmAdIKI0gqbZeHSR
4gt24zgtTaMb/bNzxM4+BiRVe3JE6n2d11HmA88C791l6TkV3Z7Azuu7nXc6B0RIJJWYybBE+DXD
5yG84p9fWEvxxle3HkCMWX/gBk2DQDvvrfbZQwG+nYWF5Icg5KnIhrMMug/mbgX0TUazq55uh7iP
Gpb0ZKXGc9eSwmAkR/XO17hR8t+NXyWgRVuIEDYW0/30oGcNLC53gomtOzy4a07TcnlQxnjG9Gxg
fBiUqRZ2ssakpyr5VhkLDhF2R0eBEvCzpipbar+Z13vdimFHTPApUIgDGKvn9eT7wqgoKvtFDuW4
BG+zk3LnKsM7VoMHJQ9yMSZQ46V9STW0hWweuUxkedHZj/a8pn4tFhRkcq4j1TKye3v7kRuvhJbL
uBnvZ82pUTogZzv023JIgzVvIfgjScI5y+S2FQ9gZ7tDqOIVl5OLlx7B9tq8n/NDDvzp6YtybCdX
+FW5SrnP7ISe5QDBgqsGpNLnMKUORfSPUX+UjaXz6n7K3PDyErV1yw1iIBXyepRYlC/uEVZ/5k30
p9RlPxBqhm1cR6Ufjfyw9iUlqFi0eSZWNnhEOkXM6ztzUNhMFH0wDaG0qNVPDCaVcubI+Ri8UxqX
wImCJoBYyeCxEFXUXdGpkmtZHpowQhdk8e0A87vbulJyMTMvkBrcGNzwGM7LBNFFaHKtcMNfA5U6
R2Nm1TvCzQIAVGC/lf3zJ+4lOTJV8KTp+yC60+VDwBfrNKlJWmXz1Y5BkIJcpsP3Ic59c89ufuzu
diq+Nl4tcFyS3L5hTUDOpEX8uQ0nQ21xDLm9StLC9ifVHIiIuj/D+jfpcoYWnau3lwVzK5P8cX0r
Ll8+ewG//gToY8g7gmgi8HeHhmhozx52zGwMN+RAUi1RE23SZPnJTpHu5nBIilMFLRsnTwrXJZiI
b2i5AwjxN7VetmuByDVwpN8bM2sBAGY5yZVEx8de/LLVHyVdwtPg1e4L0plXGnNNnqF0qp9hEpMS
71u0o5TfDK9hIW/DSfYmlfV8PYAhd7QB7wAxRSX30WkzBQJTnoPzV7EAL2xD2lw3l7j/he+saYfp
rV+cyMG0p7uulcuytBdIhLBEFCKeXMfLxibWGchBlCBbwmHSVK5SATyLwrWbyrGEVdeMxto7993O
l6iAn3oKG0DS8zjelVllnVKt79JXAik9pAGTAeDb4LfNRzxs4b70vyxBbVO3tUwAmzXwf93IwWTx
Yc9f2gwhelAefkTlKhxo6CofDEtzY/ysgoUboo78o8TMkGdclfIe2NswA3x7f8eg6BbNp3num9Qa
S9tyYn8Q1wsO37tOBsj/+VbnktZgJvYisWN7bbOZxl2RTcdW8MxQCEFsBzvuHEnqdvhZTGE4e8HT
0nXz35yEW2kVoEJLz3RVrEH5cYsEH9VpXxjmswcbXy1mGzGW5H0hKzN+3HP4OYsvZ2ByawnYZeZT
7wNrMVIaWju+MTuh30Znk04JXkfh+5k2aMzXWh3BbbDYCMMi/PlhXnbnkLZgCBBVLXoCbe+KOD9G
80q80pjgpyQwlI84e88+2vmR8OEjwNtZeW52eXpkcIXj3LZSl6ro7f+qjMxDrKkzGSRpghb0gwJO
Vsy6zv84B3WHHIjGW1BxYLnNpqEQ9SIBz1403Fb87mCMwuZVCZl4ew9mGcFqQpf82ZVcghTrKANM
dKgocURFD5j223tqFcNeL2hlNZRcwa+5M+9DIZYqKR9fHlAvnNSBvRE6RzVUpYxHTTO0FQ1FqjNL
3J9cBIZeyWPA6SikKNXEWKU1MN4QFSI/t1IlQtut9dL+ulJfmTlKlLitY+Q/Nov+cMuyB1jdo6hU
GVVOkUdrHHu+tJXxjHVRkGajCJokN+PU3QM1RSiqct00fEoXvrej/wr0bs9pcpISEz+ZcGLobePK
6Z73TBiTKhOjKlUZCZL+Qkv58ErUHPhxHQyRDBKMj2qUBxRpsNJoa0fBSNWi2VB/setqvEKmV9tp
SNQfhcQOseuSdaLZfgFbdC/god6W6R25UNbBtLsB2RMR1tSgnkwEfdKjzVj2+0WtSswb8jA3fPi7
w6k+hIVmTVoK33ScsX+emnBnpfhzxXyu5j/kwhWXHrM4+D9O7xTA2r56lc0+UCvLeUNiTWi1MD7u
xsubsAL6QSZX3VSbGxYKUdFY2Fcs8ec7IBRX958o82mcCCfeZnJ9AdhDlYCZCjOev23R+REKup3R
kFtWvCx17eVLbk4b2+7xQ9uNkGOD1Hu7ksidLXG08TskBlsDmPkzWpUCjyIMDrVkLrL6JwHYJa24
42iE0qdkcHJO06BmumKLMSmrwt+8AoTj1a+KQUM9QmPelcCmAkHBO5Eft/Gb0fCVuOS3aEACLqzu
OoyPgeSHb62VA6uxFITF70s0EBpqSlRREMSeMG3eeqITqRqOTYadjtBtyf7qxzUJjgktaNW27bpP
ay0UuMoSNnyb4bIWZCp4JgTT1IdWUE5b3PugUWRIPlfYb/9x6/bQNh89pnO8txw5HZj5AEBpEY8D
qPxww95P8di3ug+km4mlRVnfiZBP+EQSVyMj1m9OhxGnqZORP/ajFgvgPtAGatrLtzcpEB1tMZV5
PUqbAb0ZBTWK0SMUrVKntPX1Sa+vUq35Z0XcZzdXkaSsZELEa4Gg9Pk6INX+4MjxhvBtAjJvAJox
BdHcIr239ukyB1eTyy9c2GUA1/f3O5iDBCJP1G8ogK7l1yi663fqpwSNjD6hXkvOwDdpMeeVdCtH
ojnA+3tKqPmV41eTp1YuBfHfploe7zTS7tzmw21Z9EBFCByHnOSUFBft88A3RQWZxTa2UCZxXHHa
+LnW2L2x2oecUhgrkIyudRf/Q8ATuP5RKFEj3jeUx3XFtN3oude9LZ2gtGwgM27IXX/cwI6xUh2S
Pm+eJrZNeY2g3DK6SJuXR1BMfVv6/TciZAEdRyvo8VqXdkfH10dB/2a0VyQVlVh2xflwuxOiAKjj
DCsIlPxbSDX3M1+SlQsneG6CgMU6fdX2+rF5vkGwT60JVu7JWi4foo6vojFtpy979Gq+mqCCRJhz
l5xpx+zPsiCBQfsZTO02ZGKJr0hUxb69THK4Eiqp3e17Eslg4+T520B1IGKhSz5o67pKFjSIe6vg
vX6lGBTYoQa+79RinQIcjfqH/2uhy587asH9U8RqvE1BsrJL9oooQZh2pwEXtsh3LnzwK1Q05gJu
z4W26U//gU1XqljUSKSYJhooyV95s9Q0KbCCRzMGqOnEi2IXteBHmALp2zMWV4MKu3JgrdkzPdF+
+82Pm9x+8HeSx/CoXpzZFia4nCCFLPC6wSKw6BpPRCLApuagxu1pWqmpxzXMR4W783TYa1h8b30x
QrgommKJ7GCDOMqLFKwk9sh9XPovXm+LFKfLFOVseH1RwhOZJUC2c+uawkCG47B8qHQ7Bt9LSuW9
NYdXIFcx5281UhvKtHYxUGViD5gznZb5OWpCFwBEbuDmRnQPvFKttVliEyahOceT3iHgC65C6IqA
jIJWrV93NJOEbkr5HfIoDmD+XON2c1oMiHJnG1RIoiKjjmZRFnhaVkrbwRXlJs9zWKWpYYW+sEU1
1KDwTJW1STxCxOombBegDXcYeS3ka9T4d8LOH9SjmLt1V3hrnqKBmRj/HE/0aFdMlSIX1qZMyUAb
2AaJyYVXtlnzHWH2vyn1QJ+OhFyF9/zWp61+fwzHl2p+3Z1G7Y2VzN05qWxkL9sXIdwvLvjsvhQW
/Li4hOEiJCWc8X8X1bY2ADPTuOC/NgU6H2CfRdzVcSg9JhXQAldDVXIsHSGSa26OVvXI+3+F/t/n
jcsOLBZhlU/u/l/Ow/xGUsrJ4/X3L/oL5Vuw/cSHnfTGzzYStaL02ziS5vJcahGzFsZ561NqzAh9
xcjpzumaMN0m2Zq67J4ArFYWeGwgWvDckWOIhxqQfKpPsUAwcya5rzZD94n6o6YAPXbZEso0VUED
JyK8M+gosZaN5i4PWJwf/pLV0SSCICJltcTeqkk5eyhQxbXnb5MeRNkPQFpv5zYBPL7gvEdQT7zc
5dmeaVr26CSCv4BFtup2cy7t5Ik9jrBnvTEMPqeOsFwvVCWwTF2glJWS1NVdNMgK/i9G8hyZO7h4
lzpJjw/CONWg3lRxjOtIDcgs5MErlZ9U4yrDLZIRhcvrT6UdIWdOtt9NuBF9N6IWTBjsr+hnB/bm
BnEVNzb92jprr2jOIbrYX8VR57vkKfSGrrYO35Fa3l6yTzYdn+9MfNd+VJJ80c/KnuCdgLyJqxri
eRegG6ly6lAGu9yjvlgVJou7C2380AreyNLJN+HGaAG0zVmTsQlm15xHu+KVtwVW6BOsWyhefHiR
qsS53RRNe5YJevYatqQgXU3rXtcHrKdea5rf/9WVW1bo+U/b+3A/unu7Sz/E7zZCsodXRAZk6IOm
vmQ9sStZF6uaiVrpGAztJJIL2BLfG3rJFo5tFD/bck1O/7+Tn4T7TkwKyKesIvunp9BhQqrUsk6Y
DWw3LDf9uHYrLWniSH3H5LrIqUF/6PBCAYoU3eH0qBmolgobG1TcTjqjXJn4iUJ23+vi6Uw9o12g
eseIPd5vnDgkWVIiozVEdazonKOF5izjDII3sH6u99uqeejmxOMJDwTe2Osoo+ngC8gXQwLhXA20
Ph9gOH55zkZZhslX9rx7yzF9229GfpElorwtZI89Mjp8tjpJMpqIUrrpmJ8ViEm92MXXaJEfxcLM
c5jvgWhElhOn0jsTuiR8VHHkAtv3TpexCxTf8EB44oRU4TEPJ5j06111ylhbFs4efiKLmj0tRjf/
Xoa2wDvgXb9cMut4csLsUCkhjkkmz6DPegNtcShwu0icVfm2Ae499DzGyQZzPugNOvqzjg76IkxK
o3HzOcwchpSbZTZz1je7Jg7mJzvBvu/7IRZfYpxQB/U/bx564EGfgAF+M4vxK/YByIfCAx2bts2v
a+OFUuiCWMl7SAHZ8tkgRYGqwE3/EXM8wVFjd5AF1jFZlvapYpjhrolp1897GswefT65yrvR1fG1
4dcSfOJGWwRPvHtWLZphjKaD7uPRXF/DdwEgDtZsZFaDpQg38MtAKedEkQPXolzYk0Q92x5Q62o9
+MzstNpPvHLseIf/8NnmBbi/L+5PIy60Ni6SgmCPRXMhVqMYwyNl5sFjVkNq3C8J2fq+j6l0keLV
4fC6+WEyTPDtW+UqlDQI+wwtt/IOTHdQkz9ptbB/T5fu9ZUzb82t96MssnUTb0Zo/O5pJeKUDLNt
bDSXQhmCLC8FmpmpL9KzgPFm++vI+4IqfCr1hW8GqXiCc/W50cy92wDMwD8wQexBcv0S3bwMh567
+WU4hSXoJc3GG4c5vziqU2gWQH3BB44sMWmRblqr7YSa8JlpoGfX/isNwd1zQ5Qpmizu888nLZcS
gsnQttRdInBbkQtthU3U1M9TsXwVncXmbwLQ1Hxf8DSaCHJBtWbGOwRgAg9NgBz7CNTMqNO5009e
a4MTtH8HiGDtcYgcTrWMchbchOkBHtv4u0XRVVdcaiBZiGUegOddbGHVu36lUTliArNw8xcXB79L
JSN4mYC4FUuuxKCfif/94P3L9DuPLFydoDbpV8Jpk56N1cecFXTwMwq1pYGHoSO0FPs6JtFCBwPj
FN03qu49zKH21UMyVXZsPvFUGvmV7g8DvrBbab2pHSQey4DNZGpQYJslnixIuOZZWLpMGKpL59KE
6q9hbYn2TBOLFgtiJp6AkigzHPpPDyNeSWqfehpSCI/CpqEoRAw40d4dvjvN4HTpNSpvk8QJtxyt
WsDI58dYirIZFOFLl/cgw/fVqiwORGlIaBXDp/waaLDAviTyGqDEkFP0V307v7i6G8SzJ9o5pm8b
mGVUkVWgVZymwMk+WD55tCG0IaL8asD3Hx5lkag+MS26l7TG8dCGpo/oy9iHcoAr5axhtrCt+f5v
EJ2oIKc91gw2WkM1EKQ+yg/D21TKvDrgTX/s6FGFkWlo/NjKJfegHxW5KYsJj5DLBAB7xvKvWhIi
8B3wZr3zKvV9/gKBQlrhNoBSiOve7+B5HsE/SBzDRsdoCbTtuNyJAUoqlDCyH02q3e+pZAASJtrY
83N5FMGjOZ5WaE6d33tDe5Ob0pzoLeYuH+lUskkxRK5FTYzbprJGVHjcJDky/m/Xx0CqfPOtmz0j
z0FKnBm6MnZMHaaOW838ynqMy1UecrXnRRVyb/F0w142qJ7KJYQ09AYmZAtV+fsjvZeN8C0QbYD0
gB9Bq3UCTf1zv1c8rwFQr8+uOHJnbrlUlzXlGeDSuve5poU47YoseVAWJnXWpKL/XDWg28sooE/9
nP2vCMYnwbGv9SWEbw/HpbSMn/7f0jnFAAYsXITTZASW30p6VjbgSGkHEf/+hPLhJL2JMfognW68
eSMCnSCLhQb7ru/4I01Dx5NoxLlgL/+iHBcJotKJ37jzVoze0SXtt4/Gzy4wBUg7YLeMk/yTdynM
mkE/X7GSal6+XobJT8k9Qf71fZs+c/LjU05kUE4bHjjTIx6aQZEFzH4t2H3LN4MsVv65sCL0KM3B
bU4U4jBFzTx0xSm+4whqCVuB0ffT+iL88RMShJsXJt4ivQavypuZVd5ho8vJkKKuo6ayXdpERbcj
fbM4kwEV8rDZGMRKDY/7ZUoH7obJ1l58Qi5KuZLoI7rQsa0ZCrvcyYEpfXhfNgKzQG58LTIkiGVk
OtnmqrzrfnpuUuCIJS/JtEiD2V9yAk6UxyJYqPUvvsqb3vSGIZFBM1D9lWxNAnjw4gztaslKjtej
3FR/AJZftqFRzjjfS1rfKuEkut4xm7Pymfg2VDn58bdIAtijpdcq7CzKiUmidaExzVwpD47YhTzl
YNJNS+D+BEAwO6v1fEC9xKcrvLafvBjuiDElOvwUWG+G85fWGw2jL3dPHKzW6lQ5tkDa026ubFmx
RnB2guv+TjonKL7EPpTgLscdhrpCXmHS/euD4E6vj+l/4sdI4250ZEducSzcW2gr/MYP41stzLcA
ZZqeCEg7oi0qSloXsX4e/13XEHuq6h+ksdwdSG6HoGwj5V4x4rcQHSbGedku2NY+zR68ysGTDRBz
k8tW9My3+h0VUpgM6GhkssLzTNmGVNa3XbYqmnavpZV0hWbogkOd8Wz5tYzbhqzj+zpUpXyf6Pp+
jEnx1fBW2MYQt9SaT057yMyBaHBxkmAhf5v11qDY1xmQhFl6Xv0CndkmhxI/JnaGJlyQitetvM9w
VTCKmQuqaS0svznLk64OPg6CgMNwmaCT/GgHgDAN1PTB60zBjfl/kaelOjjdbUrv3n/PSEODUiy7
37zRVkh+fVthgy16MVPY094YxJ9n/TAn4bo4sQ8aMvPggINqSVZuNPY5nyc9Mde17guOHI+GdpCn
iOL0RF/UV7Y828DTYfs7/kBjqG0/OLItNl1cHO7d0jvgaFlJS/GFclnyYXunCn5gWBSDWAjcya1C
GnMBwXKSvnSHb4a8k41pgwqAcHnmBGNfoJZX/MGBKeqvIfHljZlTkFy7w4DWIRb+hUfeffN10cCp
A6+CD6d8BKxzcLdYDiV90f4iOycY0fqRv68fP1Ou450Be2kGeRYeqZYnLc2yZ6mTaFjrhYaUvqT1
ZIm6dffckPuK2evw1usy4aqTiZIPoqhVfXapRV4kvRx9i0gbvvxvdwxwjK78FvTFZtvfLc3WWRwF
QfxIs9Tp0I/hbvFP0kZa6jTFCxW89XCV2Nk481+VtteXMv6CdUtwK4JSqWQL7BvSjG0qzlWye/AF
v75V8cIPTAm2VttoavCydWU626KfoogHKjyKSSS4hlDtha+12X7D19TlFM5uEo7Ghmtl1rldviqf
2GJR5/QP1LgSkO2WZnAYTljviMV37AkUXSYTumhcw5LAxy2Wm+6ZFPd9yvJFNfwdUytb0n5lUJKI
GYpSe8X4HPDOSgibsDeBRWPZ+mcqp+xPIe+WAH6RRynGBbddCeLehbeSOSlS7en+05xAimOolehy
7Wn40kkn5N6DgolAIljzIK9gddj6LQ1JXnSRblD7yt2BWvsLiyruC7xHvY/REmwNlADkxj+PomZj
CkzIEhy62I1MJZZSGD7Y9j2o/FLxB55NTaPir2gwnr0ly+kGWms1J6Q0F6BnY3Lnh5GfVsZnTgFW
I4uEnf0iUaBN0HsscmYKbLuumBr8Xemk9PP4eCJ48twsZ565oWeAxC8KNHw6sgkaLXkqz8GDd8Nr
dw77P25ydxdn+k+B++2q2fv28btlDd1PKg6wJeotJZBYNgrQlZeQ46NPsQjUScYocTm/EHJkD0nN
CPj1Ukj2KLa55nr7do/wqs4AmvUwkENSI1Y3wy6ZPcUWO/ZKAUgJ07Lv8ZRWzvdrFggXMfivFPJk
L5iqJDQvCOU2RTqEyIfjBEEu10ldFysnmAzCMbB/cthMnVCfHoUP/PUh4WUYlBIXUbo//9TOxhO6
K7/blcUm+1HR/HUorRZMav6Ry3l/M7jpDQXc0+gen+LX6/s4S8wYUCU1u8gGFKqfr11b9g0+8+bc
anpMLtSmsH6RLJ7JsuNNAavFUN92fRYVlW8Cui1krJ+Mgvnr2JAXso7lYQvVUmUKvDdwZfgL3ku1
b9zgvVrpe1/+WbazeiB8vRJ8BSTBfeBZJ1jnT2QPWGp01w0uCJ8dtlfAbuPtLDCBNridb3FHjnYK
fxfjI3MOZVv+RDg1E5zJF264gswr1CFA4vpuE+JJpZC0tfo89Poq5rl+RHSIytH4a8gdigq6bnjX
O5W1ZTwVR7QAhp3PZEmBPAh8UAF1J9gDJLr0jmuBtCyvZNRUlV80xTDJ+9w7hPB9vtFnlX5myWdn
j6yR5fXZkwfopL/rnGIOsNED1FVeo0lR2rejEWTJViJPqFAV20F82T7LGcFEA73egFtJ5GG2s1fK
85MoUwVrqCeUym90x87Lhy81pIUotI0YpIjwwKleZ3cUDcJ86dG9Vpg68vRjCRjvbsHKl7AdCakd
Hbrb4OLGZBJkqq6fzTlmIyileMqg5z48NcaRJZOM8YjeOySJC5EFs1uK7v2DQoozQebDviPH7vSD
rnmrJXGe6WxpuW4PDL8r7hzRUgDAcFw0CdJRk+WphSE6c8NfYo7MsOmSnYmLx598y4cQDLZm8V3O
A/AixPoD5NU09bIVqSkFQJ4KmxUB45kxWfIFUX1+3S5hlmzhpbqjh6R2O3VQCFP9XUcQfUfesGeg
5WxtA8s9znhGuGyL9QBfETE1C4+e5yGRcQB1Ls2MC9ruT/rG61BpebVAMIpe5J1VnnzyJPglsarg
Q3swtCmchL/CwOAijaCQ19uBBontuG4XrjJhtloW2/HQZfAXQpT2Unyw1xRW9q+K00yP2fDAHtdP
ltXJa86pw857YlCRtEq5uGG084if6FPtq/DFZqRtXdDdjENfBJAG4NMiCnYfmWWguSlooKsvWCzr
l1Rb0sXcFvAJOEZ6ow5eiMntTqgUlGbYzANDt2YSNC4BNhcls/UQUHeGySk3JwjbWw8DAhvgVEuo
s4GYNMVxxs+lN8IM5oVmG3zapawALcrzw6iSJUQ0Um/Wafy3K0vXB1V1KZKuZtCc8hB0n9Duhqtt
NYOhmG/Fxi5uZ44by6tGy0jJI5iFQsy+372Qz6PeojYEZfXodp68riJJifZ5HW/jze4OYB3bdbe0
SVF5dI8ytpt9YeXrFZBJVc3U0Y228EZhjL4rhoGqfVwxEcP9DKscwhLmOXD2/iueWR1W6S8kRE1u
B23GXMB5VkdoDx7kiXcCMIg2Y+uncbFl30nmUzt9kaih07tAWhI11jKiQmroibcxT5kbmLsSSV0Q
BtnrDcZ5c2gsiOZmV3XOJjfUQ414tNqpzPkQOyzcDFZgJ9S5ij6ibm/LQstMs6kyKqjtcYZRXA2Z
wn9Sv8HateAK5eVj7PZ0xW80/IgYEZlPM6wt+f+px6s0TgKxWnjUJ9AHKvksYfmdLeeA3jO+SGCY
z5Eyx8l5CPrZxMBD3vBxB3Mc73rn2YUintgpyXDPdfJbe9xgE9CfPy6ZXG4gNXoBRmkTNeIipUPb
WhN5uOgRtKvjFXwKB1n5bB9bhGUSd7lo77uHcgByM/n2Fwlyk2DKmBa6OPOY7STyeaR2A7OTXxyE
Hc6fGzo6r9s9LyNxNyTIlp6XlAcqipzWnSHMDkdyQFz18RtPXjl3qgKNFUd7KfgwCvKAr/Xo/7uv
9hXvUCC0hl9j4qMYm69DnZSvUl2osjfuD5Dxz5fqdkEig0MaYMKCMM9zZu00Hkaq+Pdhlyd1Lee0
LXhUTCZkD1RM+pRNwwz24xEhROvWPFPEzCPm/lI9yLyPxz88P2zAfGYDNWnl0hgo/c38g96sh9tv
dptHr5bUIzCMuqNPYaSkmZjVfD+aPyg771GgFQkMJDeDzkUuqvkpYsOWDysJnXTXNyRKhK6eQC7u
zQciOWWW7WXrXZMF2XXSGYviGg0V3tnTPWFROynSNlDBNtLOxOe075H/a8vnZtSXUroc9bfMlQGn
CxuxCvR+BT3nZlrT6MeocqnBBM4KAtCgTAFS4rOqcnUcWiovhV5cMN9n6DrrtdLPj3iydVBIYWXC
pCnqIvGFZwhsgdOsVj2t7ExVt1PR7F8oec8h30/3wqvxP52mCpXkvcqnFBoYTyrBNC5tGOFawNg8
tOB4BRYpEU7jPuuwDqmZNkQxXdSc23/4u/UHf5F591QeP6WBW8xzoA/HH8O1F1KgaHVxScRfyF5Y
pEdGrHrIjAmEAUTtD78z5pRQZDqJWMUtr7sf914E9/qik8EJpSw9sd9n3tEPIasKzSNJIWaIJV+w
y9EQfx6OOTBxO5o7lR05XW5YR6Dq55qof8/AvkAy9WqL3LHEsyWQSpTKQWXvPWlcOf2uG9wt8Smq
gWDbezi74BXHGCMjOPZ6HuOj1LVKhX8JROENQ0hoFISAxpORDuJ2m7lhgrTTmxRgtTcOfKha4y4a
aO6vNSApfRv3l/3dkiJBMAmjdDHgA+TMb6XmO+JF/lAtdrMwjPxxmuZj8oVQuWvieCJ64bfWpCLR
+W0JSnlG/AEE/E7pJrF/KMaYzwawUdBc9wCzjoY6mJAzwn9nLlXMH8H9yYkJhdUybDW2Qj1Y2XiC
Soke0ikxPvGu2EgZ72aEK1zHlBLtvUpQ/+c+EU1pdhGe6ZkPTClOSFJ3q8UunTVLzSXY2WhwlXsv
I1O/u2Ri3n87rThxBQ2ZObkJU6N1+wIetCCIMS5MVruRCnDzPgrZkT8Zmz/Ui3dKlfZl6vIFVs19
xbRwcFatzBU9aezrG2DFFC7VltlXkBNURb3J8QOXXg5K54AijxUnT2eywUBz7JtiZQkPpIRJOPWL
n/UOdA2We+Zy3DS+18QEB95KYKK7AeISv2+YepPd9/7am7Jo73+YOcJ7vUYht+W+35IoXfUS8YTU
K0/72rk2bbZKT4stVJafFtWLycPBedJ/qu9riAz7//gw6My7/VK9Adi9lAEMISI9WSWQpn6IHVOx
D2ecgjquRNAmKGtTAdBMP9X9D2U3T+qaOHCMXqRCeMcVcnZD8APWfECj8oZRg95EzlMB/i4rUtr3
d4Sc+yP2m0vzjlgBTZlTliqK171/fRcvIsnbhF7Xv27vVJ7OroMndjiTdbN7qXQ7qIXSLsSDF23+
EIgrk38LTwaL64bHGdV3gt5Snr/hMxNhd74vEWctarPyHaSdiL54tf4Miu5bqrih6FjXlFEFmPuw
koE5GHnNr484Et8Cv8UTIoTsaoinFdBykIH+hXtzAAbKlppRieWQ5L2uEq0Igwfy/vboJVWZY6YL
exw9NhxXiLpBbDN52lMJ/BgTDczpZk7BfE8xP/X5DyHJxpnppwFiPqUWqIlm+IXgmzV2AzijpMXO
2dT0iog6IciTOKTQLiCQKiXU4J8CmuzJ9qmjEnmTLfCTSa1c5cPxejTDc3ZFw6EmAd7VqD9yJEHf
3YMfi2J8W0StlJY+lHlzlgLu3Dltt8BQEBEGTC0WQNqQ4DalgtXWqJ/zozDu152HAqpD0CTKSbhD
gZHOlh7yfe4qdUHcN9iJzrv2QCi8n1JGtKrwVUD0Lv/PRQXypv8NPuT9WgyFY1qQrZ1D5ABq94XQ
Mwp1Na/mIcporBg2lOTEe2KjXXAUwAE+tYbssDJgA5cFnstIy9wLXs0T220fjOTNjZiWtxdFxoxs
A7nR5sSn7fVJncSJ1/Gygjqu0HxTen8tj6ENxtEtN5t9ZjOKX0LQ5lFovT+24kssg+kaZlVT0XWN
fHWq4+Q1A0AG1SVbXcmzObVgR+2OTdwIpFZrGabeV8UD9n8wL7OSDRieTRIzzklVjNWBIJTkDJPf
xBAWzepAee5Ok3UQPqaKJ1UlyuCJhSX4iyP5RVY/IZov+DCJbvZy1ryeeett1D51aGRn1JPX9XLU
MwM/l/Gkd2Dyf/IyyNFrUupoC9c2J5DWMxuSbcLTbowHqVaX/0maT36CTBQ+mqAV9dzdwrfmuqUk
MjTUHoVHqsVIyKAMhlCy+Y0hXNid/tgbe6ysZ2eWWay+mwu/PYchoiY4pv6lp6pC3o5zOeHifDh0
7mzM57AwgCFQkMmXj5lJJt2whpRT0c/Kbcks0vqMF3O4RlSbl1JOn3B1LY79+BwvZsIPN4Oppp/6
TJE3w+zbHjSSz/kF79BuhXgr02MexEBn+m3z5s3yssX0VBfjNGVU1JgDXV8pIB73qK0pj9u/9HtB
ubwikfFSaZlmTITITQZIdBjMlMQ6dqgH894mvGgqFMfn24RYcSL/9xXTmhqbld6CgCJ3N08TUmZM
gQPMtrsNR3DFMunF0u/a1qXAbyDrdPiUsN1bX2/FCuLApyAjEm5cQK/qj5PIvr/W9VNi3BwaLYnn
M9sp6LIP0ZwNsnzeoMIT2Q3JbfamHdNSNW9Lxpg3ufsIahcQmV95u9+/b7Elj3DXleC3E22SRkAg
4AUpdAJumAX3Rz/Qg7aER9NEpkFwukZ/MX87A94+s2Auj59GfbPSBOd58LrumOTC/VyfwxWF97XC
sXJjSXDjsBfM3e91J1E7ZbcPOGRGZjHWKOVg9pdBqFZQ1TMutleULtLK9eo8O6CA77uHpGI12OpM
Cl1n1HLKFr25QTaQT7YHiQaUycGjBrara1Hp1kCx3vUeNY7p62mjSM3I6b/9ehCFfacwNJ7FxpLu
+b+jnxIVSNZFQegnleIAPFCos6j5kcNG+kCAZa8k8rGxFBsDbHh+y2He5anG5FESkwsn+IBt+V2p
ZINDJEV/Q4KPbz+UMbr9w5KXUNaJ/k8I/bCoUOwaTk3x+vMfY99rT4P8SQwP7vQLHhFeSzYCGWpW
1TriP5yf9lum2LSBUUMQhCKJu8OWjV850nxJsNwFJtqnW57zQ942oHhGMGlXfIQE3yMagh/n6VbB
OzisPlJwMVLZ8Y73BPpe9k62GgWS4FT8IOvHp2cWaRIU7SJDFPwqaAUTbMzDJ0FxTxFYAqPZAChp
Txs7JdXIZndQsAo76h+KhtOjy8n/pSxutQYTCPVP0ya73BFSakYhTfdFqJRR1LyaeJg/5qBLrkcN
JcDBJHvfkuTZXtsVqzkODhfAMQd9Rd5QRbI8HNdr9vb1YTW3GjTQQvu0TTincSGN7BE6lGfVcBlL
/nT/iKHXjlH/ijxElu57Sblq0ewrFZVaABTR1DRslAsaNNdRYpFku8fTGMXLUravwvf5jL84iRD6
yniuCezk55vVyFrL0PUiMg8ifmA/D37simEy7Uk6aL8OFYlYL5oTRz2076km6anI59eTSPcv0DZ2
ZzLIOIYRpG8gsrj/f8GfaUEO1dlUvSO8/PBp8rl2ruYNWTigZjgQTOcdSC97SHahKikf9kh3T6aW
ExYF21CDSMUzmU8EJFHh+C3x5wuRCBlUFDtp4dh1vidjiZfcyH6EzukARMV1xn7wu4nB/rr9Twdv
yDMYa0AxHxfCYZ+W6kzCR5sTvA95luhcrttKsWWcV3si1m7tRgB4V71ARRU1FQkRsPcVWXJdBAbH
KUHdz366yG1krazkwB0wGWqrS+I1+jsVXMbeLWjsi/2ajrR+Fv6glimbbVcLAXHQbPQ/O+Bd1DWg
oUVoalRqg4HaW6xYp+NnQ+Z9l5hy07t6ZUKAZ5u8fp2RS7iwjmZa8IOZxtPICFC+3z/j42Zh2I8c
gDFDMMF6NOx6NuF9zqgfbKsVAG+kdiJDMJWGptYqFn9gYa4WDiNJJzjmkCkbzD9hGhscAu5heyD9
9oCFmKJ7bHXmPDGHXm/p4ibwNcDpLqhrPJFOUnjikkctUJevRa89VwoyrTztCWM2x/CSVzzfo7Hj
7/AlMV5+58aVCKvL3lhIsy7y9DN0pqEShLXhxNVPlkN/axWUkJ85XRYU+lfLCfEyjj3dyFeQRrim
oHDOGbL6NWs9ltLM9bWee8WCIVxSTK3oeDY6VNVVeHyD9kSWPnFlxfaX0afK86vn88gNroroF/R+
lmtPgZyV3C4ZA1cpHT/KcTKItfPdi/l8ig8pyMEbXflHXXPhLmiBF0Aze96zJU8r3aXEc2g2Kv/m
nsy4/d0KLhLb2DqAyoqgnvzkG9SDP5Vo2QW8Xb4oLWtSNSZIoXLoL0Wc8QiQJ1XxffzSN59xgHVm
kwBAqnqKSfm73XXCJrSYMl/SvYChhiCzIvC2ypYmJh/lYofJvuirUHBluWJl0ac3VldhIXk0sv/Y
pgm6HzmXQfPWXE07mW2+YduZ19ePWwyVkyL19L8YgZsdIS2jSjiSdqyHjoIzwA8oXBIdDztru6Iv
NgoA/XOBY5Eso9JxjSPHAODWwQ6VQIdBK7MBiQf8RqFUMCgJdkM9itLasjco5JeJrCn66adCwt6S
AhX7rt31DGnBHMkZGHQHmz10X/U5qI+18w+Ot5aW17x/3gZyAp9WciPF7BG5n64HVldE+E7P2m7d
1Rjmr8ouAoZQ/1LibZ1irCTxFlZPcyqXhkAVkQMrOqcZbhkOKS9GCSe9iGkJ9Xt3qfI773Tcx5qA
BqV9AbE8c2I/3BMhNPMYDQDX6XgQUlYUoePosaN6nzTvio2ShY3ty6OOWbj7LtE9DVAB3S/mZ+JL
OVFONrRykvBcDEDzAZ7w6Dkq0gkLuP5n7XO9HlPPV4x8Yq63DsBIb3lLsWya7G0P7syhQK/SaRGV
xHTlyLYDkXXT5RQinXKUJkd+Tx5waAOLJ/HJ26ndkdjQc7KHd43HLhkMRUIdJW/sWMI5rxrmtCYH
Ga+qRkLngaUYbIEJXinRN+Gsf6aupz4T+O91wYQ6RifnC65Q2QIyEi32TvfR4IWrrRAp3yi/ZUhF
FTMW7g33EGr7y+M30BvRXCFP96TkVcs/a95FevF37S134xmicVEbZXDxUs9bI4mKBHiQ5vrULW0y
1h1A+f9BFVB1eQPbnxwCkozgVGDCu9/p2ZDPExI7QmmQePExriKpQPw1nApYBKKaixmgMLrYpa0P
xy1ehnB71ccc4DXnVEXmhDytMrghphK5RFIDiI0saAAMa7qHdOKB+vew1tfkHS6VF+vIfBJcylrk
fxeKfNXoIExCVRqsMZTcy4+bEiZj4ILMr7Vbr4FMkUGz0ljOWpSpTq1QuV1M1+MmYC7VCwudmB49
fHiFsAJoo7WAltQZ8Z64dLc4exSp6igmvjXkHpEcZ5gBtoqEoVMTnY40RDcSlxhOI5LJxOEmclJ3
u3VXutbIdiP+Y/2CQV3sV20D3xRwfMcj8JOEVuIJtACKnyH3QckaxWnjisg5E7SiuETaQRA/dDip
tmOZomk6OuS87jQVnVVh+He4cmKXQmbCGjuiTxwmKMAAkpAF68RSRQPzXxKV7CVixdpTx+Ylln8+
4X3kLs3fC/n6zjWeOxXGwmCsB04nOuM17KMX5Y+SMSCSR9IorABw+rXFCnyhHdQ9vdPB8iWhCPYK
wkQ8I540JrAF6bUn/9CY2fKSbOwg3bsaAWCPeO6Oh4CJJSJABClkB6EKINBEOAR4GkWTxnkdMr8H
ktGoOO5llZTqjcS8LU9snMHzcHOPMYB11JS9nbwFNC/efFweQebrRBVLDBJv3a5ZT6/LEQKhAo45
YfUbu8GmQueBp1y4FysZ2R2p/BtEz2snrhEMJXoJ9sHibcEd0gRdMmIMDWQMoKer+dplE9pwFF+N
OEJFLmlHuT8pOwfIrmq8tgFcsiWzV2QLsh0bcsbKPC256D1HB2HNRjC3cEyPV/5OVWYYZzR10H8K
+BY/LPEZYzpGybiVMvusR2a9SFm4CruO4aJ5l+AcPR94mCgcC46PHuvGR4EkYYsTysNHYtpXEsy7
+cHkys3F2YqpzK2sqoN1DYviuNB0jDr909Ka5RORQ0QrlRhGcJR/pNE7x8qlR6qGUTq2/5ttGhoW
77DfZ/q9GVm8+7wFqPLFVOrv916AnMI9MyJFQ3p8F9/SFEW+gG/CW5r6rYU1J9W2sbcf1i87igD5
cOXOLRleajavjy34wFsalqLWmAkXUvzMciv+MJXOFCvfd0LCewqe5gOXlO3I5g3KQHuK4ZbXZk6E
uFdb8E5Oq4QgquRko5rDf8LziCINjTodpuo9mCxzSVy+6qMNjDV7qXRMzWGFhp2ppvbbsfz8U09J
K1ZazWfcCRzBm6ke5pfMo9/PT5e5ua/rACyO2LheDJl8nos0LrY7vKvi/VvdYNK9SUgkQlJJAZ40
+GaWLPYRz7fZWjpvlTj8D2GxTRgWHPUPZEcWvoISy63j3IXc8OmAFq2m644/wh4CJpwOZyTTMzmD
wViKK6o0+zoHhUNlOV7KzzN8W/xVGebAsZJ7qqAHcjFkv8kIczvnknka+KoBMMCZhvAXoUyAc/sl
jusz4+3TDPPSESm0+PPCzFBQSmvkDoARMAePaKkC95E2pxfL6YQFeRpCnVIP8BIjdY8wW3FMqjum
Dhp6xNMkUDgiKaOhxhe3YTxglN0u/eTLEnZj77mh9EdYtnU8Mo6S5oIwrjA15V1WJSdAHb6eu0In
iOGRu8a2i7XH1oJVDr+bQMZJ9R4RiSq1AXhEs398i+zIMUKecCuCKut944vNPxc+PPjrNmqrs5xi
QYVI4mDbnUfIUSY+RXEEeCaYCloxhzhGJUoMB/7N6jrVBxJseZ0Zhhr4vObhorUYA99q2CBvftdN
wMHgw7N2AIYQid8vOVQWgz7LipoGYocZ7w0OgoLz7oPuT38NpiJXsEqjigNw3YnzCFRK6uH9UM9S
cA9aFx299tdW6U91BWspGLDVor3ck1GFAxlwuuna39IgDlSRh9ewEhrfte+rOdmrapPupUJAqfo+
lguyNA1p4BLJSQ+tVS5riDlT6I0+agJw8XlP14/LpZkNA3lLjFzPG+GZDTMY7bmh7wr/XIKjU6oB
++RHmvUbF8x3kvyc2+x6U6ZBfCdauOFVFOAi3qm4Nw9Co83f2/RvR2qM+2RjkbGlShJBGb0DgbyK
CQCemTLSZTzjeEkVEVzKbDff2KEiHmfYX/SBEoYeAmrCmq7RFk6mOMPEXvK3MeWQGpzjEEjFDYIu
UuW8M9j1Z7EfYUtUg5JeRdEGT8S0R8ba1EECnJV5NKgfh/z+UlkNwGQKvkB9kiG8YMvkoZrbZzYd
UHrv780P63+x2YgD7HIwwRY5mbEZUyfg9jRUK3grg5NpX5Vl5I1HQiVLUmx55rwxF5M4D23G/nox
3geY9mOUrsobIxENLwvw+uqXIxHELweYmA8zkjGaR6WJzxSCu5YYKj5lmyne6DQChUgCfq9Sv+w5
BNfisTYFY8qCYvf3LQxyiiAGomwD+BVIpkhcVGLeBudCLDTQ7nx7J4igy/PD2d9H18v01aJiD0da
A00li7k1Xh1USv8NK5tlOnCzTzgSvZIAv8ggZ35EJ6V5tjME3T3DxRLZUQH4XG5MyMhWFGFsRgDD
hEfEbs8nLJPEMOec6MNOsvB2KxY87zTatHa+HCGHyg+rBVlPVFGySSjHIyJ5rLgaDPZUCSi0MTAV
JxFHYD3XdWWSRyqLlTtGxpFn0rKe5SqHX7sD6FOIWKE1E12OaEfhPqyIlt50Kp2Pho3hDOzd9Whe
QT3GDWJ/iSGDyNzEj7j2YBFFZfpOnP9xAy6dywag11vbE3O/xREeKGhvjjLBev89rSO1AaXYFubu
9w3YG81dUDptx5NGPfpVmzixhntGQ8Zl5mPklExOgMLnTj6wNPHGA/CNSwtR51VvzFb5O0YD2LXY
PBuA2U/SBgp+Rzi6dfTkDKifW7SSzQj3JefUAAnzTkypaGO1yj5L61uH8lnxc96RUtEKm3rFMnvh
ciWPX/szWs3rZDJUrsIxBcSwRLpz67U9PNSrpL8eKcBpmR0ljwMzOSlFLXCW0RXbxsiIhupC5Wbl
+hM/nyNxGOMjBJo+++Vb2csBsdkb3glsCAjsDPJKiZPQdnjKs45suKC+ahQpTxx42+HWxRm2QISr
jqsn1GB17GhzsVrtxMqVKlXVoO58A7kHXuzwn72JyIvfjagpbXcwagbkOhYZpl8N+wP0hZMIWXcF
W7kp5fKv2HauIvlhFt+KnmiV7Y81FLodSQwhVT8hvfLusn3KIRIptEoReR6JwoczbSRwsd/jTBgb
yZeTN9W+dGKXKcZzxwPDEZllJUjYUWjfVMCq4rTO/1nK+t2SxutP7OmEfPzuCSxfUSyCOlq2N4SX
+It3mHE91cEuytZC0PIJUuVfNov1a77CWpots6tXp7J3efS+XcbbAi3oaDJTpaGKKXW12YJ2ar+E
5CP+N+UZ9rRMAmfJhLgp/YTWDWM7LUGOmE90cniKE3Sq3SwVYuQpgBeNjaDkoSPS4YOY3CqTNoGl
E+J3LFXQF8l6YjiP5SIpS6hqALqJqmzoQAAwalpXRe6+C0vayl2P36oDQGki743Jh5+1mkqt3bvc
NAmHi2U0kivyululwQgUf7KyLnTo6ubSnNEwNZAaxpdwkRS7w5WLn6osJxp6MHVJqjNTHKd9ovI7
Xjsuw3oUyeQfgGiwfXr1b57WkdMlOzagt3k6jqGoiLU5yl7ZRpWeuA9dfln+DTkNSx0YKgTJKIcW
KWJh3e7va0FYMZVK2+86QX4kTKWl/l4tkOtmrk7TetyKcUNMWnY56tkuFopNn7AKgiD3R4OpH63P
S0FTGWYDOr3n/OerrqQka5lU8Rjmvz6w8g2FxOFQgziOdvdG9Suhk5cQB0r+ETRO7fABPQW5JbbZ
/88imO8rFkJaolsZ4UESzpmXkz3SrEQYR99E8Nx+xzKwqKeWapXIqrIJ4vIYrAK6o5sRlM1+WSC5
nCLlbwZY2cKSNRcooDtNhtxsCJpF2UEJGLa6DuO1aGg2VoJcWg0s3l+2+4NOwTgQMLOCr4fYw/gE
hP2BUCqEOIM5iDgbTHhq5LhfVunE+pWtDxTHiQG+rBnojk93eDWMtRS9AGAmkgseKSF7z2CTgKz+
FiqtBOGDGL/H6dUusdDQ/v2nOHmQVMhtP3iAhtR7mQXSImB+Pji3zrPTaCeZIwsl1SMlzbDakIOR
bkD5aw+p5oJnt0nC27MK5Dzp4Mb/cvxy6vvG6Pwq9ouxmfj9gTaeE/QXQbkDRWdLfFbZAYhtfSG2
/K0Sy1jqKyM8bIGchKcgkVuDu9zHpKGXFwdWMwXM7iXVpZoy5vBai34C2tWJzmAc4BNshF0Bf4Ju
h++lpZ7V9pi6t+gpuSMyxGI8e+kfzwFzCDKnCPirK1ND8/gkJjdwiHgBc09uFcMXpUSlX3e3gdrG
YFA+7N4WilJdrMTQq9UshnlbR5GiBAJjneO2/52lJNHCn1S+2a7aEUjEnJwyCW1UJWkmOPFfOVkd
B/0X1sF8KSedm+1XxpXhBxxc4tzqNUe/ORt+Apozwp6bOQIhYs2+TOMamGsuyrSU0QDr5m5vJVia
xIJXYfZhHFQP33ETGpQp4p2KqVIzOlOOWAW/yWCvO4ckBf51yNvaYuMr9t6M3Ecq068FsISVS6Pr
G2GJEe4ehegr1Bktw9ktbCc2cL8ITXycWR0N1huLMLjKDypICT1bBNaCiz5IfZ1b0qNdrIzqX3yF
vs8JYbdCyWdlWEy5uIoJsZI5230ehf60c1n/ArBqDhAIFHZZK0N4clCPH5TUKFlbFGM5kGZ9CkUp
ClnsH1w5VcrZ3+cV66ao/4xUnzvrs1wHjlSojFkzVObCF6ZAYh3OV5QWkl+gsOHRIJ3XUShx0zQX
vxKuSOHELzA3RCnb6md8l+Hfggznkw5oxWu/OmQSo292yovITgVgD4yxndA1A+0/O9J0/4uhtsw4
8r8C07AyOD91WLc5TE5Y1ZWlWTIeK0+56sK1Zxp+zkipJd8KXBSNDTZSgsiG8ITPe2pQrlJRII/A
5Obnn3JzseErOIURCIZbKbckUeeLCPQL3VTXNa8UAqPM3gcnTGzuzOZNRstSICyWzOGedLkrAxsx
kd97B83HWKmGHkvj4RRV31VzKKKpw0l5pm40S3VRRTIQCr6bT6tOCtHbhacNbVV2+dIwnbbXCk4B
aM6ETgBs22sTdrPPRF9tozuJucQvL5VFBlczUFsBncVaptjiT7f+JdHkr6WJ1qqUTS7SzhZntysT
VB4WaouzGiRoCcEANcJDy4xJW3M8TqnyfVokl0pau/FmFC8fS4r9UZhMn62ay/67vqvVTWMx7Qdg
Zthc2hjPNXZiQKIISuV8K/bTPypvAU1H+d+nNbXVOy7C4LtPedoAnlb2MfnNQ+uRKw2cc+OEnV/L
xTMn4aJIw6TdlNE3qWQH78sS5tZ6WIsJzFgvETr1JNGrfLW6d6VGWIFU8+IWetvki/Q4JIlnMtdy
XW5aNkKC5PY2cX9lfYO7FRnar02/VAosl6KqyVpVRq5paFTlrJ6wZyL7v9o/YdduUHbVjl3uj9mZ
KM5/L3GrqUVz09DghzqdWEec5rYUm/OqU3YPw48eAKzNChwQ4gzPm+iHzlnYh9L+CUdgjfPQWie3
LuwKBpXwODQhhXKZB/Wjfh5hp4R9CNQcUYxd/CIwYFmEIdO52bDN6mwQT/O5Y+AbvdZc1Rfp45VV
ksG6INpTwbG+ZXXnivsUnJa57N1hdJqmCbP4doMnJVNP5Sdmt/U7dckrAWJDK6hEbDXjF1t7iixg
TU+N9D+60MtSAfiOaPpbk8wFyHo/GR863IDzjN3Hd1lXAfmCF246EBfqY5G81WqxbHyyeOphKWIg
koDrtPii4XTlw5+3l1wMRH35P/g+cB4jBFszP4C9YOi8xcENvXyCWwWuizr+dQR1eyvX1/qHZe+P
yk1F8D1A+TOZmmcsBrF698L6xXZsC1t4X0zjr6rUe/Nh4+xSMe6OqsZJGrtO3jKLpJ3hFSJ8rlG3
gEdtTFhzti2UlcLOyULOQd6bqsUC84eq/8oTt+A2JXzR5O4rTCb/FtYoocsKI/uhrFe5f4yQ3qN3
wA9Z2sjGLIsTKi4QjukSNs/WRzcmrmldFUGqz1tIMlglYsgY4XypaXnyxVusbs9ADBkqgkNZ+Yqd
8nU6YGGDTFvf8p7SBWowhz2j82ewVSH7DRfGInzbFxGXrik+PVTzYLgvu1d2lb7+1gmt0atA4PuH
G9ZPzwOcK+0YS/f1Do4MlgwaFWDb5I9S8Oqb04zniPUlzj5iCJ0pi2+RESVak2LvT6pc2Fc8SeNa
dKY7vCJADFNwODsS/v+T7T1MedlHFAHdKuPqNgK5j3XQv7fmDD5rFnx/3b+08AJefu5D13oBzlb8
LzcX/z7VCfZ1qYny9zgmo2ZUNHvufv4Ws1V3NTg/OSgiFYqxEH2jlFjZuWY34xMESQDFaBCr3doI
zG1/NQi/O4fp/SnIQfPs+bhc/pZXqyHSLYt2Pui9+ziO3gteyCVb7dYBamZWhQaWwQrfFe/IbmOP
8nf6bD5F6HQv2QKsdn1W2ZgBkYH3Ad2PhzYOYBX75KyHHyWFACh8Vz4YWGr5DBnXreirBqd59gVa
vPzxtgJxUGvYSa/z87+l6XMQ9Yx9vpRpllML4N3T8nbN6HAb57JSRIS8643xVaqVv1bkJr32Ygnp
Fu8KQ0jNeUSe0cnrRX8kd7MBpPus8MNog6Z3xCizX94yKfo7rMh/OgwJ+nM53mSyN/yp3GBLSX1h
go8e/4rKDvPRx/QYX6sWDVe5VAbkzxj3JyrqBzD3Ukr+hy5ebRVcu+L35UF8PE7BL2Ln3TXpC9/X
Y5RdQEBlcplDwT0YTKZ60xdqEMMNel2kHSBKvmcGUe5NW81Y3hf1dt+QYEhdqlVYc/SielJjfBXZ
xfX+AnH+VRK8/s+ITB7TzwSFf7Kc4r70aRrr2TEaJLSBuOgD0pgbH1Ou6m99+DJnSK06bF7gYWH7
uTJ36BtU5sGvLIhEXyEZLywWobt+JwSKahUhvASOslyHHSFtL8bnmkqW0U+uDgALnLYDV52pl6rP
TAj6CeG5M9D4EQML617evishwgP8nBeVyD7owTC1Xm33QQSyUXGa1JpFSw6a9ik0VweqNHQ9yJYw
AQSJUX/wfCsdUrx77R3IWS3RfrYXnPiHFiTUeZLsfKBnQwtv3cVdUurKU8UKYrlZsH920pBkCfNm
OmJ3lpLyIuouWq6SQ38lR3UXMk7rSLpU/2zuHLuIRM2S7lbR+3D+8KVd1qDq3X7bkrPoCfLGUFMM
+WHIBOgozhaL4/Wekld3CClRBZPuYU1sD2/tAxIRdlsr9GfX8kvFuL9UZFd1SsdprLf8C0z5U4oM
shMScCnGmGSZLN2FDz1GDYGEQy1N6uvBOQ/qSoJKvu+LPcRr6GefMPtyDU1ypBQqlfjiVqGuY+rT
sFxsqZwzkW4IIWLWqIfM53mNTtgS3oQbxR7nuQTFMuHbrBa7Xigl5N9xkatgSGs9Hd/hvY2DakB0
sfoocdDOgVqZ/bCFcPBSeuvToKYnTtnUecepOlwZUCef3Yun57nwrxvuV1AO6y+ZdhTaT9Y7O6vP
pv0rtwJfGMjXMaRtJtSRLSCmbWLAy6iLdX9Zefkgv0dmFbzpyq9OdkGLtFn6qp9OOcefanMCjwiM
cEGvZHQAxHLO1ykY8/soSdFXlC0I4YnFftSEprrCo7aYBXzZHluM9loeJh6Nysp/Ilk29/IXfOaf
Bgi054Xp1FnDB9WOgY5G4w28u6cqyP+t3aNoAB9JwlNsUZbLXzPnyj8yLc0I2RyAQ/i7x0/WD6Fm
XkIlNWy/7UX1s+CH1qD1/+/+ronua2D3nsFz9EJDWarNaIgNRQsBld53eB2Bm9j+pnFG8eNlAf38
Os/1ZXGpfmGCr4sxnR5EpM9LnB6Krs1SreBmO5LE+q529HzHmjSOG7ZAxED1vfHfqtEGlYN1ExpO
E5q58LxcKvOhHb6Yu5/Fc88Gowz2Yt2V4HHmt6WZrbcKTIvDtE3qsFLUbBQgEuqJUyXk4b11EOdJ
724Wdo4ZfJsJUKkSvyVp62CL3Hrm47qeq0/Y+dqvz6dAv+QOgRn0luap82LWSkbTfgH+0q6DSXCT
A3WTBYYEgSfR7JEXkqs3dsIdTsjieQthfDqUbMB+rH5bSirioVp7HEH58/rjSWsLCuoKT5dpW1Yj
TTm11T6IZvP9aeVSB1nzm0GfFBsp/PqIXS6i2utjoyUAhL2Q/9qICPxwmvd4cdEbghVcjEgY+Zcw
TQQcg4YwpKx9doDwDxTaaLRMJ8eOAWdK6CeIckXbGr7xL4KUETeHFVMd2Mdr2Cm2f1Z3LdzbrQ3U
oVmQUUbkBu2ILJIozlc2B04yjDxSPwCmT5N9K22EUHyShfYqpyYjWQvmWkU8IbOSdGNzLZpZEMx/
L8kohaMbPeAWJXKxRZpYmaBODx3YY7MFSiwvGVonR90KTIR8sjJ8ko6q2zbDCBF0OFHUK9YEMYnc
6U2+nI4ZykndzSBQG5qRHLJxvRoxjzOkdJzds6nbHxKWLkzSckv2JVwGSMDyUnrSRxUAmJHb77K+
yI9qRPRn0qdnl0BiwljzwwCnR1htbLpwiXUUAnlyex2+YflhXfMyQCaRnx3Z4qH2++ZkTEeNe/wU
I5bgM62SaJh0EntJrKDLFdzhJ2xM7HwL0oZ3HrOGGdhfLzx9NJhbkoQF7jrYqAGFi5CYrwak0xNx
+Yh/Y8HYW+wspCsMeCPNnT2U1MvHcqTA7D6tcIot27rvTTSyDCPyr0jC/hBW7ELynQKIrocZ+mS1
3vX6lkqwDn+CJ5TNJc06s4vqbtbuPggV9yMWTrS2nCRH+KtaJiQvhk7jcWFevwNyl/1Kas8S38e2
2HpaD4qZGz7zAomNXXquD6mAmH0kMQ36kcHOYwXmZL8mZnrZB5Z0D6naumdVj7l3g5vGxvs53Vx8
zGhWUFILCGS7Sk5W4cIkczzFLB6SgEBUKRQOoyOc1yCC8m2u6a8eJAX3f8nAYH4xNGQ/iLRxrZ4C
T37AeUrzm8FKpoCeOt9BIT5/1FrWe05PgieJSQGw2BoziQ/814aFEYbkPEXj8Nh9L646O48a1wYw
OZ75LLAMP+d9v5cparkdC7xmMGgXTlOF2KdXt5C6AeU2Dhtk86XcAP2JLs4RGeiqOFNzzACZcSPx
qgeHpz6ZRfT96Nesy5bsp03jv4z7HdanVvq7qDiMPrVc2sq2LDiArkJrwGb9xOTXrAak5a6ZpoSb
YxoFjoUj+W088Gc+pXaz9qbjRngQA2u3xoNhjQG2fN93BQJDNeZEznr3h9wR0iE65hRR9Bku4zF2
jgyWaDDD7QU2yf9G2XsHGWludM8a8GKX1bM1vO+NADBUurfJ7anRKZ3GApHiGk5OxvnAFarPpGSd
prLVn3EztCsQFGAEm4CTuFErsPhb97Fnrjae18sjwP/DN4Vw3Jr9HP+LXb+OwKrhrpCmeSh+KCu4
tFeRzi67hzE4FGXLOcFDCF5X+DWZsNVezCLfU3jsLWXo0Q3L8/JqDUcT3xITEJvop2fqDFxDCNll
KHsLvy7jiSQUdKvUhbbH2VVHM7Xnk3CT1JBZHMRyCioHw8FLixDp0F5Tvdz8DU7lgvdm/GH0Qi5g
/pSLYHbmvlXQiedoGv/daVGLy/QuP8LRe61Q4XnkZW+cUNpiU1Ac55Cqe5NcGqMvmJgmMfqcGMm2
u9dTuG/3gD1IIWbkD3jQyjQPCsh8laNZGctd+nPlkDT9sNdOYpkYjziHBllhlucqteAzRaXhylD1
1whqhtELSKLyoTiyg0a2hmE2zO/SlZqyHj7p4lDcNxaJ65WCPk1NvDiBgP4R8omcHkJvnGnl0D16
9S8CpRGcyhl0VlGFUz/trWtqCcsNRDItTOve/JC8qQ4Qz9KyFVLH4xlsbzRvSA3eQ4X7Lu7oG7eo
YUupkY/S5WsV5OZrK+i7upEA7LrR6Fcft+vif1n0hnTsrpmvEGps0Wzor2Y8dVU81yn2kwXBNOy4
/cEHRU6QxQHRKb0UQo1kuAyMchMv8RIC+fdwSuM1NYSwBYY/d8Pmu8psiHIRJPMK2mV2L9GSbyW0
n8cyZum1gltlGLR1PwfGxBaJJYIg4O2xxhpgdv/7jsoe4DnetrvMUo6w0NrzkNAqaA5R0zfBXZNR
Ms/31rM4IxUMkmvJpTIwVl+Rb55zr+LrgyBfmr/1Iqq3yCPmajUieJxcCDQEjXF2JM+tn6TMNZNl
YJiJD3HWDNUUd8kvRNua4/rNrpsCAjwJtQSea1IKC4brXARgQdR0sfAikpPDywuXn9BOFLo7D2tY
driNrJ9lwDHd/s4e2VDM7H3hNRTkq+P84PkqMCeoseA8v6Blj95ad2i4xCwBMQSf47PC4hDljiy3
Onp92weH9R1PA57ZV6d0e8vQFxpM+FcU/xV4pF0mbweCBjYKWjFrpANC4ndC4S3NYTjSOLU/uOG7
LQNLoEG3SO8x0CJ26oTM4Ex826uSXuhh+y9Is5wurrBUABBCLcrZRRbzwKKy1CpYGMhbBMMt4wo0
rn/lBfp+narDKpgVV2ea4UaRBmB0SyqXGZI2drVzgkxADCrgCHhyDYucRwyOwpXxtwru6RTKahdT
Qjzh37Wu9XL/49MFSA68a7unLVxildRhBwfop/Bz08kWRkh/0W8EWOn0Rm85gLC0XfFt7b5pAweB
abEvCuZiopZd+qrGu+omNI/zIl1tPIsy3PG80EIkxOac0Ch5IiVyTNhFFW/oFzqK2ucYute9ecm3
uUU4yPURK3vL55f7XP7uHgWK4T9cHSOHfp4f25vVlgqwT9DR6aZUsSCw0iCIoNEQN7z19VIaCy/z
tCBRR5m+189kSyhJnugYRjalspxqAuoL11YBPO6c0ZjUPa85JdpLctfjTSsMNMPmLF142lLJMHMK
jP5DgBn8OJIxD0naLV0ovSOWMUkxkuqoxQWSF3yeQf1hIgSR9p7qsLMwWGoLsD1C5o745pO3Iy/J
iTHkBO1QuUWoTygoKeUJNh9RC9wRunnGvNv2agPlyPyRr8ib6r7k9M45L8Uiiw6lQUP6VsmxS8aZ
lE1ntIwK+RNCVqh3ErscEG0bXT1C5F5SdlHtQZhVH6AkesdX4Hk4Zlmr2eRmMC5mbi24kylolb7O
kghKt0vzy9HmVJz0HQsnuyQxnMrP2yrSnztF58VXFb5KG3nVo7dqmpZCbek8sKHR6icYbXT6e2zz
Wu/KP/KYKumybONXuY8sKKo0bK37MEZZIwhEWYOeewY4nMvKmPWKxX6hdycJrAsg+RKP0iXxRVfz
k2eoJG8yP0d7gdDJ/S6GeRKt5Qww1EOnkVAXdcyGH2u+VypkadiVsvw0Hmlda2Gywh6zX0vS1c9f
FBMMDAYRJ/uDTw+XckwrIw57tNVAydMnWhnj9tgyZCBk0OuUbwcvrbbxJtAz0TZvqENGgM2udlxy
A94O9B2mJeZwPgfpt283vEDQJJ1yatmdPP9hSUltGZ7hqnLi64VQlXuop2+X/08zS2uRwf+LX1DC
iRAnjUmIBy3SLBRPc2O5HnVeBPG8Y8SKN6xHg2SCPOaHTZVA1FazLbU5jejSxnv2YX9zm/YvWupx
w18uSwv3b0Hd04Utt4+FzZdmia2zn+BuTtsfbyHw00g0RxxS+MZ5c4E7Qyft/IsZz4cufUyJ7Ynq
GIhk/O38gD7GgilUbdzbYZx1DrzMiLwBzScSoptPVfoesNcRQxtMaoCY2suvDaqxBHzaYb8FuCxw
PrBuzddBDg+TEw5JX/Q1LNbJCEQYa4Vw6Ng+EJFdHoeOlnflJ7O1KXPL6JtWqOnt7Idf7fGmMRoi
S/Wb0eHJL9zTr8FQf5IeutMn9SFUIewEcYEOpDmQnIfK4VhkIRqKTW9BGZSLx1yjB4CztQmoSfOS
X1iU+itGTAHWJiRpOs5GcUcEIodd6TKNNCWHEn52y1NmKz7vW/wweEXjC9z5YVjChQghmrlZ6jR/
DX7Ji8sVw2KQcCelXvKi35V2t9amgaxl2jmehgHUR8LSpAN30IPMt5+EB5b4PP6IGHMz/IyiCsCv
d96c2XBs17Bfol/mykFUFrS+Ny639RFiV7bFzLNW+/oUkIaAont5nhjlQLuF4GJic1/8NsOYvf0U
NhOOlFTnajFyyeSSo4DUqoBLKUvMAxFYYK5WPFMv7EfP/SJoorp47pJRSGJkEXOuiThWR2+4S8Do
DnauN7oJvY/7W3iEr0OESqY+8sDMRJ7ydvucfpRnqjPWogqylcoEq8bEJwn4AHd2d3yHiHc9ptm+
8QdVEMhSwsmIQWe2FduaHXHKj14VKvIBEWCkMhgyM646kWxitgrNurZo0I4BiCUJQLocTzWJHgnO
ZzBTKUDnBwEEPlKQ5iGFl48XTBhlaoMlO0rGuhswaGpQKNrcnoQ8e87Ua1TvTUgWGlLF0LfJbHTs
QdIcAnPH56/8xss3cafR8AySBRoD6Wd+vFX8cmUNDX1MnMPdDVhR0ZV8FF941Q5Iwd1jQy3w5AQq
gv+CIGrgmFMM5HRYGInzKcr/PEaJ80CsDg51Sc4C5buYmmyOz86pNNqIi3nl2lgGfaU1ySZzp7Ml
LeIQK1uU89NLHF8uNRSW493dySM7TTPrKK9Jfp8q2xAOby467fIopGpACzZYGId0mlckCCiClr9O
nNPm4bruagNPuj6oVbbo8v3wfXMR3Anc5S9xqMmu0IRdE21Ia3yGk+5QazPLskVl+6RT8NU9BeWj
emzV4aTBDZ1Dvt7JahVgGp2hMSLRm7VahRYVFU/2eNEDVVQajLk5WaxvBIaUI6hzL9+yxqB0PYcL
PMlwJ/yZ/0NbaNrodqj51xKmDjHSFoz4btW4X/TDAmoRLuLd5I4OwGz+5PZ8ACmBi8V0Vq9qNWVB
d5U391emxKjKWJDNTBG5+INJBIH1QtWiapfPXHjD4bkQEc1e0BqrndVrjXrw9kzlpOIUWeBmMvyp
FYPFInr4V09ErbD7GISDzkLYf7+vyElJtDyjIEk0qJ5kUrrGFZupjJCTG2DCeAul3GB3R732UV11
lbxMEdhyFZy1Q1QaTO0eniSSp8oAsXuaGA5TOePfLf6trk/lVVBLZ7t5f4FeDiwBYgoKpMgQHjVO
zHWJvRd0LucRiLd6walm7OQxCW5CF8VcFV0kIooRvlSCcFAuI8OeBLaqQUsVA24Q5u/Bn8LfYLdO
t4denjmSVFd0rKKYwHTzwXHpJtV9Ovb8o/zpKEkWCF+cafs99EMLS/CSS9Eg5XXIggaUsPkNNMw0
zW3AVRaAilmj3xYEJmuCcpmWsHNsqBcmfGKqObgRVLElPgEKBEAyqwMI9Vz8bNqzthyPLThL1QI+
jlmBgQ9WKc40SmDyN7TBoxivUGJgsKF052FQV0ZvTNdbsU2md0Yz4zwlNDT41PxazuUhyuex0bSN
v2dJbKoRIZetEHHJJXGLPCOvm7WVmwDsNz/HARmjPKb20Ts5xuuXQNzHfSAr+D2fvCDaSfVPwXn1
ax2NKPDnr7rRY2S+HHFNwRfRPa9sJPIPJ75dv/ToYOjaWDIAlm42Pqvh7hd3CD5eSPTsZdjyAq/M
2Ts9wfT2A1n7GBskYRerKF+6wC2riAcqWshuuwW3njCIayD4zJ28L7Ixv/OkzfQJp6CmsGFQNrtI
vVH6du7brfOjq20UG971OYKqAgGp60KQ5hpoqUI8fJK4njOX+UIgEuwjHZVkOoRiosowPn2Zc0jm
vGuQLSQA2eFs9RRKtwlpDFQkSacRWuUN18d4EInaeFFtwjM9vIcndfrqUn4QN2nEZIo95Thz67jd
WjGZbtuKtwvPkbjdNBKeF4XW4JRn71ltMqPB2rj8RM5gY55RsuNdLjNm41alvF+pkx0JFRuoKDBx
SwwJp5teCH6edkHwrdFCvIoXrO0iQ5Z6W1D3vKWx9MbyIq3NieavkKoeRecshRS9FBrCRtPQ4CcZ
j0VmyPSolIS9zdJL8LcwTTJRt0TdXR7tmr4rnyNp3pDILH82Co9LZc+0DSb/IRjjXC7KcUrZr637
iylnh0jdDDUNqXBTdNckc50znFBfcQQVCiqvHQuurEkV0vOjiUhzCG2DmVcaxdHmcz9ewLwmaqgx
6ong5KoD6WCuLKIQZQH2mpGivEdQpzB1ASJrDx4kyOHlLCkPYl3v/CU2oCJsKz90eoaMeNXCsuUm
POssdModXHuIv1AsrU2xYBgIpW5c1lzTvImRLZCYq40Gjnp3XJiv4un/0VDLUkc14i4CKKcAYy+1
EBL8GiCConOjb+ffcZSYmvLf1HpuY7YKAnR/Noq0vxGoIabAY46FAoAtuWOA1h0he33x2agVrKcU
mMKM3FnBQc75RCU5TxXwvYVHdJYZqEWwRsuil8zovEtVul2Xx2Zs722WO3UMvNSTVNTqtDjNWKit
CCyHi1sDN3HBgNVRa6QD/p9AMCV9kFdLcfQbpBxeD+suXs8dzyd0GYNtmN01KQIMkSL03XSHM25D
GdPHp4IgCKJ7RpXntkZiDsZle6dwdYPRFf0I4n9v9c0o2XIPW7z0C3lsXLneg4/bPyoKihf4Im29
R0BOTllsLLXPtpFmgpoO3kiE6Vhvf2aOxa/t6Dh2ERNWYYJ3TThWvqydp/Mb0BN70+bR0+kXWhiA
AyD8sFbkSeXz+W0VkuR/OX4IHy/9ChPYcr27BWE08iUEUFtFvkQ/m+Yfd0CbBRXjR9aVYkNj4JTf
4N7enopsTUq1WnAF0t/qQK4qCna/urjXGsJM7A2uOL30YTyXvMBZfiPr4wx9A3w7r8vR2UzG/Phk
oPSZjqOQTX0bKl7fbBN5cbr0vBVnaWNx7TTev3wjXiqkh6vSMHzVQD8k+YxwpxzUxNFqxDpGYbBD
9ZqkDQBmhT9907IR35GcQHAtZDjKRl5b0EKDF+zzmDo3Bn7/VmALl1cyy49GX1fOpAf+3FmkGX5a
etKrEou8xruXi9MIFX/6k3Q59YKQgNrsCjkESaQJC0xW1o8utV0JR3yv+K+7B4rLwKAKmuPcf03k
nGaoyNCE+pLVfnkzxI+I2ZH6lWqgopXEfUfSrpWuvRGOduiDDDHc+33wz7w2SURGIortOU5zzAnB
LYJ7YRRbRIsBpnhtchpzq7eMw2M0Ndg+IcWvGDP0fUs6Zl8pgaSdC8vTX6axhzQUk2ADhdt57MGU
RnnG8hu/J00YMYBFRwBZNjzB4JMq6wz/DiXl4SjRUHRr9I9EOs6P0o8TYFRkNhPGlOylW5bmeXva
eXAqCdv6jzy7bkvAENg2xYt9qqhp+CMlgSgu5DT4ZszH814tpg8Vmxz0nQTc2Hd1BY0Z6M7szWVQ
HuzK9OZi4CELkr3GwndiN5RbAIIND5Li1WkuAVq+E+s8qv7aYwdk6U/Y5Ese27up4OQSStF0ftGH
KVZIOauhtg9ro4LbQXgIi4KdaL9AwlOd/yp2g62LidkfcrqYc/mwsKfoP5y5FFU5Z00WKVtIYNdg
VrlQ/sIS0IQl/q7Fzdbos1R04nYIaAoFnW0ca3jqzvNCGACMQwZ4KIhX6fhxpix40y9Zfhb1+OgS
Te27N4hP0fiH5xcZBPq2tBFIEu97AZ0Q1LiWHLhK0YsTX5XZqBqPntDuvbf5tYy0bvCxJ+dNzR5C
tzeVfGU/sfHzRD7Qi8mPw/v9YHRtr9GG/DrLOZlyVzVwKWANW5/DKWzSWzGC1n/aA7My9uEPXtoS
XcW64O1vP3t5aK7HamNlYjsDgpkut3oO5QxNjNTpas25Kdqn0kAFDozQvwfpvGEbKVs9Ym2YeouX
dyDN/atuPaWnY6MXOdXIK8IlKeMehX65txj0SjywFkUfLP5sbU9W62Z0H0UT54/VPD3hymVtQ2xy
gDq28OHiAvaFzBmHQxZwOS1YkeATEKXRbWrL4vOZ3EogR8qR1NdsjJ0MJAl6BikxMDFiRMJyaNpH
Gqba2IzGj+RpeczRLXpLxoFPvltMpRkTmE5xSk9BDKGnNcxPS+nTCcYRQ4qC2ch6880XTCIA0TiQ
PyfZAjQpTydImant4a3dpy35rkaFZ563Au5BDgeLafuEInXzAm9Ex4WjZtDKeMOY50GRbxudLDe6
q7i+6xqJb2r227tVUdordD+QCuXVnCd9ymgD0gc+OfhVlkBM0joAqfUBxBUfCPa8c8NBJ7gAIqdV
Fhc1ek6pBiOk8kx9yPczAVS6fHCX81hWjloGfkOYgK510Td0Rj3DuzKm1Ia91KW64Dil49l+6Jpr
GDATk8s0AyIJ3LHFKRdfSKl5p7tYCPRm2S6NXpEvC3/2oEjDi2EyY2inp78a4dO306ggIhF/5LJ7
zteeciP0F710Thf1DHJC0OelSC1UMMnMJadHKBgiaMG70JtiOWcavGWlLmGNQTNfXyAN2tElwsZJ
Da2sggXEN7ImXsMnsEwmwjNV61MdaMDHKWYQ/QJ7/IOI8RknGtcKKolvWPN292KpAr/jys/IZXcg
PGXSFi0tdf2r5kzUOgZXYVpbshSZYqx4uAE9b7FIrZE8zxc+UwoYjLLJ87S6PgakFJzsarUR5+1K
86CszuMU90/1KuIqJX4xr6qRjcdve7+zeA0ECYzKb92ovPyRV3KuM/lGJyuFK3KAh1Jx5ub3X4d0
gNLd++S9p2frDFXsXTUucjDzbkvVpWqDgJadPF2Z6u5rln5hf4Q7MRdmfzUOzZR/NGKdpZdjywr8
Xt36w1Tgeo4sNw+Z90t5dRWxlaEMww6ewwWHVzQGxvKe6JK5w6egS6e05iR4VxlIeqTcljSRQyXY
WwXCSfgkF1IwRWyOcd26h+qtGcu63Im7ceN4arpALVsZC9W3ZdOOEg7rDHwnNpj63I1JPxYISKqY
SWh6z8vdxeZWU6VnpcIc2/8p1HjfqAEauNIo3y0U0OImJZTqwYJBzEavIt2rY85BoL9mXf/biACl
hjxrfmMZeehZ/7juSoaqjqm47/kW1VOGmMbXxfhXXwbZQWe5isK8rbBzsQslLf/+en23xAFoSgxw
fSj0Gtj7yS+ITweSvgzJGleDr3Zxdi0gL9FQP3xaEjm9kwbv65Ya6Bp0f+86ph0NC538nhIZx9ds
aR15FHQ32GtgYtHw35M+MsCcN1lwt0AgXzTOMHFh2iPu0jZyutcJtrZdX+XocTPJOqwSnGzdYeSc
m4UO/ZylIlrVQXA1WRDZW/j5mQIYVVsFuWQTeWq+6Nmo3p/IizzqY0AW7JZ6RugdqM0xYE6gFwkW
dGwtmjRQg40pWkpIY2dy2zY/ZJTDGpO2EUxkY1PoEgj115AcegeBzZ/o7nk9i4gBe55rz96yKTO0
keCxvyAdahG9PeofLYGsw4E9iqYK8MS7owsNhRnMHCyIc6V77sngHIUp1Bvqcd4zY5mLQhux8d6F
ciypiHAtk9O5VTAsAL7enMFg+K5kZ7DzighIloaXZ9QH5AH+DcIjbOWrltvJHSAl/EV2+CzXfV8b
PJ97KeZbaWlbNXNGbl8BaIzO5xPj5Ry/esLoC01ZJK3QDsHQ1r37gB3/0nAtO3BQgZ6CtVFZTdcP
PNJZ0kjHcUQj2kf10y/Ue9PLA7dJFOFxNwp2f6lAJ2u52apX5dCCJQMaA5WWwGCqA6rUISj70Jah
QmAfQ+bn8UjUykeqjQrrk5vwHiJLjeZskXZAmZWXgOle7B2JdF1EG8aIuxlCtxu0/56nkvtya00j
5fks92mL/WxQCQ8xnnM26VRm1uVmjBGHjIWF5uHNCHsTpaBgLd0/Ug55WdMnS/6bbRIbULvXB/hx
FV5WfkfmmHSUOg0F4gfSZTJ2lQNPLUV6bL6OtfwCeEF9vd5dUVZrxfIm8DSjYaVgKvUGSSGnOmQ1
kat7AVWDiLWZz3AQ8iuoc8zSzYB2hIKVgJUq5gND8T+TUND7CF02nPo8YcK6fQST4RKvMa8SYH1Q
XZrQ294qn2loYoWP5FJSd0/ucPscyARk+3+5/bw6WllcMlhN24hQ++QI2y1+g+km3sExBAY50YTO
qxAOBqiJk29rvxnWNAY4iLEdkdSPH28PFlf+gwG1k4G7cpZWwQAMlBD5N5BXamXVz27eT2sdKoxI
tL3p3gf0hrIU5lwFfBRy4SQVnU047nmkq5sjHwTx0UBkDrELOxHg3aJmK4+6ubCZQPmJhVFVbFA9
moW558HHyxw6NqWTV3wiHrnnH8TZt8Hfo0q+AvyV2W58rly50nVt0K2GR/nx3vZiGaRiZyAGTQeI
AZn7iMZeqveCYuq8uyjoiL3zSkJCY7VTYQT9LIxu4OdiDryQ5GyJaQv4RlEcS9+YKTdUMSDR3w2c
1/7dV+O742GTrnmPl9iotuLijpq1pmA4vLH0jvPk/xusOSKdwLSxGUxxZ3vISjBbkPjSwUvOAY9d
XIZLe+nZ1hla8/sPoQEvdavvaK1c1DH7O/lyu6uVrEcHEfcc+JXYDk3Bg/mobRafcdJLag+I5Y9/
KakppXLCijQ8eXJwZCa2rFyl/d2lpHRb6seHB1IzM1ppnEUP8svgmVQ/gIzBxQc2EPibRcCx9kfF
k0AsFnUJV2mrbiXvoL84ULxWrWhGBJ/oHb4M9FSal3WveK1Q+ZTVgguplfJi9QVd4lyyxIeT7veZ
lRnLnEzsIPirewtYXL0xoUf1Y254TW4APZA9HPWEV/U5h3WPRN7ELSpm+0q4a36Et50HDqHH49qk
DFTR9TFxxKV7joUljW3Pwz6Dc8bZqx9FxgO9ZOIG5m4iH3YrB8+FmD+qQ5e6VM0NxZCN8LqHWL6j
G7aXFJHIRFsOtFSxm9UmB7YYRi7CN0TPmLYUu4OSR/MFTnrYunmvrgeq4O2ie9PQI+VXzBBf7i9x
TgkHecO6PZaknS1kLCls6kji86wIPs7oe+DG6sfxdzjs+Kv27ZBh5jD5vW9bJz45zS5HAoT4YSvm
88S6RROnh/qYqgJAqq3kDOg/oQbxTiB970Abph4jH23rqGzpPoyLLCTnd3A4/zcNmNGhrOmJ5rP8
1LxsdZVGxbdmBXEfa1TwcSSr/pfanfK6FG43hx8hMFwQ4XpjR7KyweMeob62fvwzWQfZFYQwsFKz
kol3vFCeblOkEj9x+JHYkqZW+U6r4OfJT1yy/fv/Ol/zgTsGUya6J3aRhQuQHHy6ia0gYzA4ZyPW
GHFkDSQbpPM/E0k9e43B1mWcwIKOKjdODomuuMq15TugprubCIMPKMuCy9gZxNbOuI4LGZWwWSZO
+pOh9iYr2Iqh+MigwO5f5zdNuUjXqGbUNt7ETxB0djXFlP0OfvzGLukoFkoDIELFlP/mQy0lspKm
IsNlmG5k1EMg6Okaxm9xrf5BThC6I/aL942g2zKgtdBTkilFR8SyRq8F6ZsU/s8GdsPsHZhLB0pd
upePz7sMoEmBhBk4dnUYlaZP+ocqvdIzHOKhx+Y8zZelqkKDlW3bZ7gsGT5AGAEyWksoFrYY1oAE
VCK3CLq0e//YLqU7AMkcuE6Wzcs4xoq4pUnx3t1YssSOo5jRM7iiFwxl6rut4MyxwtXpSFyjQl3W
Tp5VfovI/As1G+qSXFhiZ/lKD7zlutdPUi1oyPsHHe0TPYJOrrNcxIASVDgDN/oFAHUBtBSOn3IP
Qa3LvHNN6/KMIyMCDmp1Ax27Ho+QePjJGNL/7zkOYi6xXPFjRVFjdnGWJyKf2BFETlgZI+78TeBs
VxYJaeP81fWEeHybag5SO8/DoGHaAatz6IWTE375b4byjbA+bh+bk9MDrAvaUYEGai9BLdOfjngf
C/9ckC0tpV+O6UyG5QEmyMxe5Ct/3yRf8wyerNJJQLRLqAv3ln7BCpXf7Q+QTKI4i/3R3r/B7NSP
cPbBFYIb5Kg8pIGwJxj2R+JjrL0gXV1ij5tSjDMkHcSDElE4x2zCl2BCRIpkQiX4rDM75blgz06T
V3cJ8uctaw+ECwILAT9ialIjl+qmEPQRP66RAbOQuqjTAx6WMpjzdwie3T4iHwOjUqYFW/nUE/+w
3nLVdNPJFBIdRScxYKFXxnQU6XZ4ihBMuzbfMfDB0yDPd4jeeAQnaRMSN5P24ytAGVeON++Dcx3+
p1jRJc/t/RRtVQirvpfYkqu81IUyTe7jP4W27pl92V3Lk5RxthwQOfaQFwQKyGGDPMr4WOrXsD/D
tsiVv4JYjvkKPSfSTV7iIdgV5Y4O9yj79A+xKRVhv7+84g+CIzbqJ5rYOxQ3WfFIuEBmhASShxo4
m6FRrcsBqnGad8XOxyLrFWdizaFCA01eS2GtHv/fJ6J8/QKp2dqaGZCKuQ6Bsaj5fM0gXxbL/7Kg
wb2A0W9FGWhpBS2GlJLI15y706IjDhUzzi7JGIrtG1t6Ax/0RMyVRYYDAR7SagykNubGSgiWTS+G
2+DbxLunpEQJoIiSbZuOGTYGbk9xJnohlFQ/AbQGAXWGA4iMKmxLQ7b2h13heUtQNMnHBAao4lNM
WN79Ezp10Pv/q64nl12C1IKW3cKkiYRAw526pWi6yWtwI4ILthGktMRJNUgYBYzZLUI1zIjWAUH/
IZ5kg7XQ0SdlC1S7PfwTRYX54a4jW1XANNaUf0E59ihMGXGbqOeE9O+do6lNFC/GMh9n+4vxNpIb
jShoc0lDul3aLJChVCE86H8FjnO/ksDKKiiS2rSG5EsI63Uval0+4XgL0RftMhiTSMVadilJl0J2
OHRu1dxUKKabWCTIfUFYiupki11FyEEI81JxX0z/JEFWJdUtk9bneCcAnkbIJBh4tGfPUctlAEs2
y7oxVmtMh/1ORBtCJECZAmYpAnASHuyD3Jw8qw7SQXwlH3/dvyC89QYjRs0KSVKp1FGWJokUnctv
Hb5jjUqzsBMjkLkzR/4bo5oJE1wOMsWrDK+2hD/9Dv1h45iGYS2B+kSFy/466DpJKE0lwEaDNJLf
7vbavBVnQPcdTa6FY4cPdSwKFvd6QBSS6HBaJbCehjBqnL3Lh8zPvbklpaJ047IvUPLDQplpJvu5
LWToFApLp36MH8nEKsRvG5uhx6nONy2Vt6F5kfJHEqvMZ4GF8UEzJA2tqOT70FQA7yFs0IC9FxKJ
iS8+xu5oZcAW2DCF099DEnQdgiHu7JJ7MvHp7/Tp1TZLzN1B3ljwkVYQ8yL7GHmm5cg6xOGqXCJa
5IWTARP9OHlPidEdzkXX3+BkOUKaUCXkpHlPnPXFT5TLlMDxPhoKUd0vYA75j9dQqlLZvD/FrAnh
E++C/Pk1hue+ivkjSzkDQl1bGE3mYJ/JlfLsJNiYyAwMMg1hGPqZWCc8owY6YgLoG2q4y02BXJi+
JlNkiJwafcmXNi4gghGPd/qozhdI7yHufuHKpDveO2fsSsbq4Rsy+eWzhuXKT9FJnEt+/fnV/sD9
evOCM3E/R+ViQTrQ7n+EEdzNv7TJVaRIqX/SQJxmGuwMRYQJx/CPjmxQmo1ncVfIsdsufTAkpn8y
dXt8RF+EYKB6d8qXcirfJL3kVA8YEYtYSQ1O44OQwudVY0ovTNFGWoQ8T3nS7dmOLpBWpQrQS3ew
GGmSKxvLrrvdwe1FnyyLhbDDDXde8yHk4zkklbFxZ84FPr1yOjudH80KyqbUQ+AYBa5/Go59P/8L
23gIgCqxNhvp+RUvUauy1qvMAQoIvdEshxbrg6jQ+hetKilZCM3hCDvEV4fDhCMl+JCda0ScO8bo
F+WCH7VCx9RZe/CSiECuGvUCwE1KZM2MzfsqtodVKurXNYTwKtS6hJe/BMAtUGacE5v1ro3nUPxF
PkQlDt7vV4d0sk/wKad6m6KD/dUvO6pwT8vQDE34ZUwtoNX68aMAfZSEIWjGJWL/Xpu3nV70dfJE
UsmwLUR5AcjK0ofXhVWYtHHZr+oJUzBrLRo59HBiEHwRZ+tiBIP2MaQfW8oK7I+HGNTCHcPP0G+W
qABEnu9XsW+FMSIG1UhRXHKt/RokQWeL0GNGRkJQhMYXVPpyS6t2uyrPvoQkcwyzt/Q7PU8bQAIN
/lm+ct80pHJqR92GMEc8IuMH+8W3ur8v80NyQ8V5IKtCkD8EfVGigJm0yasUEB3A6VYPrgiBf3xV
oU1UdMhHO3N1iwpkZfFNEPHbcr3T4a2nX6/6Trwn66cqS/HuGaWYy30okHw7/6hYfXjcOmFUwyWs
+zqDsuHF3iI3QcwTI5d8W7+2s2o=
`protect end_protected
