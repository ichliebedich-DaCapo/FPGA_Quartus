-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lOQtkmIXv63w7h0Ig/9/dETChMlX/J7ls610ral7rC4IUu8eAKULnO7VYTHm/kzIjjyY8h1HNotA
4i6MAqTYcepHXEmypDhvuoqsE0GzubcRozbsULoJ1QJKrAxLcgJB3cOsxaYlaIm32llNnDrkoCJu
WRIjubSG7udvgpOnwBb5kPMqQkgwavbe4RyDp7h30SOKoJc0tEbZAP7SpxykzXNcaHmOZYxoFR5t
04j9lN8hxCM/3f07WfxnHHmwf2rMQ9e47BchfXwBB7S6JtdKjQMV8xUrLJzjis/5J7Q0522PBQUO
2Hg16TjxWGazYovKssP+141sbOK/D6mONUM8+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6160)
`protect data_block
5acS9ic9wXqr5MLl/KIG6OTjWad5yNbdec7rd5z492Pd2JrPCLw56EOcz1b6DfMnPrCultKPIcWy
f7/54UyqpM8faosXlLvbtdQQrdAVU/8Nlj3rcUuJmsr4ADtZ0LXmUq5gUhmUPUM88OcwhhP1MMSk
21BFuZGdvvoKS9CdE3NTCGzzJyRcF7RgHxVsa0sXxEyUZb6/HKtBQWHyBqzRgBvksRuyGwk/WbBF
4C5QtfaQyismbLxN2Srrur1hN0RMfUvti4OP/D54fCH0n58zPL6Hh813ocK9/VWj18iyGxchE+m1
Oi4OZ69EZEgkqCDaQIj2ZVJV2tzr+/X13o7UbYCOSVhWMhRLqQ16CNixRIzzIw9joDezp0+IS9m5
4SanFCC5F+KO412aJZHCkCxsL+HIPg602A+X9mxCk6KR6Vjp7KDb2lrb2Ppn7ocjfrgwcQ53q4VF
QQueSnLPM2ZDWo/vr8YP/BDvH8B6/dYiPsaSA8AXFL58768ictL+la5nQh+TwSph2ukM4l1FIljU
9aTfEi2OuvtxrQRIb9x/5G5DZ+MhcT1ZX25NWt+uKZ7GSqJjHBDNJI/SL1wGmykBnoxleYMMvoPF
Y6g/jb5mDe/ka2QBZYhigTVHaj4ghxzhUAfcqq/uUNuC0lzYMAmxmkjQSBGiOi4oqQvpCQJt/iGN
Ekx4CTTBa/9rASBRCw4k/QC78ld1CRw4+/YPu5sl4zmZbMPn/m4iybxsbjDHIYzZy9w8FjsrBHEv
h61mh2h6VXe3yV+9HWErroKs7P7ecNA13TTn9oVolQkKCAkzDH6eYzjimVpDh/alL9b4970n/Na9
LWSMnCHgU2j6o6V+IGO1ldwDZs5MUndo3S7y7RmbNMpjbC2+OC4+avT+lANsq7U8/b7JthGl3Bwi
NjXrfHyNSXcJ3rCX8HUEeLNNYuga3NXabtoIPrATOgAHVeEO0D1+wq0CtG3eFOuodZZykaDTcLe9
rrOFAzOYIWWwxN0dzYXUtUXP9FS76OrnbRRe9lEjL2FQo0Bd9BMAw4FnhJOHUH0S2x5r9CXq7L4P
ualwMzEJ86fzAhfmVKtu7FjwT4scCuU9iVuU1GTYjVqdETkeVaF+GqBZAx8Pgyotdf3BFC7fuXe2
DWNFQZywP2mRfE0Go++fGhTHXDO8U27VeDt01/uIv2Rv/KErc+gApX3zElerXKTVGOwb8XE6OInA
0IIWgWfovu8vm5++I05TLdAuf+ZyqL1WiDJPRCsSQiqSuShWku4Ir5TuBoCsH636qemIGCHiOyP1
sLG+pF83sgog0H4wz9FrCrxKGWBRz/sOZyLHLOJmx6VQuDCScMjrBp7lKrKtREoic3dohREcJ+Zx
LwKqK6lrhSoO/3LgHjPkJRznkz7ZtVYYy+yrI/10J8DuQncVzd7dyXbsjze0Xy2mJLvABbt34lDR
+8wx2/01/CQ751VQ7SNj2j6x7SBfbM6rsDB0EMhe3Qjo8Zcb+UJGiVlRO17SfBs/H4razr7IYRes
QKFJhnJgPidC9Ucm5lwJ2NTtWM/mZHanD74jfSP5Dryi33udlybaUfXatfCG1+xqyjbxYk9LRPMg
QmXAeApLOxk3R5DpG5XVL5v44erhav7VWcVFM/Ftm7Rxaaj4kChHPwS6EWrF0PM/A5CXOMYEEbFc
0Zd21fYcCuN9ervDev/ivw+X8iI9CeJWUn2NEZ+At6Nu5rJ00GaiWf+NxtdNL5RbPBxeqznkbcfm
yQzTGjvbOfxt6ZPNy5kMdDmhxIGWNxTpUhrX5Dz5/21BwucJTIs634w1uaFvvri7fMiqeVolTL2u
H+heXL11s8FKKMzymmThn4CC8cFajqPxaoYl3YL2Wat8no1o7R6dMES9I/KjBv7tIWz2BOX10jvW
ss2GRplErHuvjS7njZhqKspzeylB+N1MMLzxPES+byhXRJpUlXtVRCzNLWo3oodR4uiTC9fgM7P7
8V4+OA6OcK3U2CEtyWyYT64QAuYo9neO4rSzv+0+lGjxvwk2CGvO7RK5YSLxxR0KazGQGSo5Qq5Q
dokLhRSbnsMNtjw5PZOPf4/+56wWpQDRDpB3Hfys5WtAfppxgmZNZ4faQMnZl/3sOv+XVzE5IP2W
PAaYOu8/a8Pb1ai9G5zJno1K7+WLVAIpCtDyoM9K60+32kRvZI0XpdEUe6Nz5pxUzdSYueS4gw5j
GmV/SGJlXriOMk9nNPzgSds43oXyYalwhmZNyHNShpM8p84pNHLiEOvQhriXGOxvkhuyT1tMlLcv
kFbDQEmcn3UIF1fvIA948IO42qJiARKrd7tnW7MC4fqePQBspTcmaAskcum7hEoRTWBUniXECaji
wqZph27C8Canl5LfTADj4jtEXOdkxd7RDAiL/3UDwbCzBwk+N3DenkwdxcaLcCJRY2u5p2/DezsN
aTmaw/cIvMyHPX0781izMCd4Zc02QYUmKxpHpVuIKXQ61u0WzpIYQ/oOyVbLRu2lnRWwco1uNQVu
35z3+7xiQBCXuXI+QPgXHAn9qNpWtFaD/9kjhGpVlVsehJWOqmyYPegEfh7YsiyBpGR0WkBCDOWi
RNb1y+oqJmQpSDeZGEDvTEwLnr+Ci7mQlk0ZEtDePW49Z6LSKYloEtALkhCxxRFnuFU72c6Bls2/
Gu955E/WO/pf7gutwjS5Daj1RXy8tore+tXx2gTxPu8WZGuIjwBP0rmnjH91QSP1Z6HTMFwuui7m
+liRIXYQpD9piajdfI9SOd2nz8kaAcFbN39gsVAPHYmy8G1hqbdymq5hA9bJiqPGFKlHfnQBiAsN
qBXEliqEKO+G7EHDJtuFPo7dn9sAJetv0HjOwjhxodhk234Q5oFfG0bBsdguetujVaWzK963f5ja
NBKKkiTsnmjgarz5DCUUz1WtyREdrQ5IneXgHpQWu5/QICATP6d9sJ95Ez5ZjFGeBdkmFlrsGbnQ
SpJnm4GYGoDmxK5wZNRAO8Z+M0A5NNAHv2yM7Iqh0oBouyVAQKMg+a8BG5GmBQZZ4/vuSU5dzdgf
3jYwHINgrnviaPJvpY8Uxto9bDhsxxqihs6KhQyB1B27lvcIVR7g75YY4724VsJYY1QGS6jlxxah
/AufTnUK9iFW3w5JIAMnHkXawMkXR3VEmTdawefNWQoMOjIq3yu9yTniTmMORA8g3P90ytocoWjx
Ad30d+f8ni7YpLlHtoI/XB00+DyWmZOSMCSirgrAzykvQLoymlvcqg/MRKocrM0i/xWz2D2KAMEM
uUiq81YAiMF47WovtBQpRUagCy73p2t6XuDhO3fEYmAsKOwpFgcQW0A8y3xalDNEb0v2YGg3gxIR
C3HRAmUmImdZbqWhUWXn+ki0yu3/5Av+oiULBgBcjYl7I25mPIgaq8xyVJtouNZyMcBnzjczpQSH
qFElzOwgiEzJ1FHLiGnGNBWoLDc9O/K/Xot/hErQOw1a5Ihn57RrIBAKNYHq/IBC0BWDtGUk9yXQ
FpGUguFwFJjAPd/q6pDG4QXwKPYSsekC4+zM0i/Yc7XnXVL6BVzYiOXwnqPBVAyvzrZp2BXFE+5p
yvi3i1rebczYGF0XjEUbXkI0i/LfXbkFR8HRISPsU0ujUSSIY0frgyMXTLbn2U8qq9b1ZcbW09fm
vObQR+sB4yq2N+gD0DE5w0DfPk+wXZpKCcqw/5ixjYEdj0t70Ky+1j4JBdfiCM4N9aHkr/XB3GEY
g+LDoAK1ZANq84kyQWi9WuMRA2lBcZ/t/ReYpGrm6yavHbqrBMdYSDdZopSAW0YtKsUQqJMjl4gW
eJZctUblK6NV1uADYhzBqabbA4BZfKZkhdYj+d0g4ENdK5pNN8EsPUL92lZe0iP9gOdN7/9WYmdb
vb76KWHMBh3WpoB/YvF7xwYE7epbfHYQpLek/uvivyMPVG/r5yzFptQyst2NNQ7ecSbnQ6+kGI6z
kLQTFOA5MO9vlGKSwx2hIsBYxoc17EKwsetZI3d6FMF0BydrVGkFZJOnxMzO7oFeBNlrx3P8LUS3
ABZcjOOioJliXv9Kx4FCFzyG5whJkhgXBQ9dZvhjt6b+qi7RQt78+l2PaWVZvnQ4aeaY3zf3NOjh
q7a8hrOH0egWU4RbgEo8lmNg0yXqjtpqRytcR1vRyeh1qAoLZkM2jpGz2Eta8AkLVmKe0FMv1h8G
e3vgSxpDD+oGFPFRZZmTt2VeZsz2m19cNnkcD/B0uVLw7JuJHDCwhg4hIsJra3S0zAL8J5xtcsxO
dR/b/ECFQxUAzEi0T2jqKnbOqTxw4rjc0gG2Ee4NXeJL+MPO7nhe8ZQQQEzcq1jIsIWaya2t9VTL
mmTjO/OS+dH3p/qowZargN1dWJn1S9/q5ktknj2CMBflwxXldDBtrHh1sGgF0Sd5gglni4hMe9aw
9Dst5YIn3Wy1RI4u5c9BmrbPnxYewkC4sm42s3SZ7WaKTDJSOeQc55FFF8zyqPGIxcrZFdqIS+ck
6xCbOxvg+ZnZFqAmUTEhySzLmshoBRiBs94XBSt3/rws/55fWib4dboau1R9XGRdAnkFUt/KiIRh
oR6tjR4QXs4dTvxKxxfgH8mMIpWPwW2FUosBs8J2KPBM/NiM+nB+UkSrfPeCNPlnU0dv2RPCHC9e
fCrTI2Jc2fJnGGKaxiBnFCy6bI/bYsA0KEH6NNctcPzvfwZkt+D8vbLrehoe9fnmOm5zPSyMOYSt
KzDYJCpGrKX6UerdxecPnD+GzEZaxxqVy90cvEezjTqQN038cn/smh0RtAxN7aCqrNW3jCU23Mjy
LgpqITb16a5SinYoiJodIYZsY6XNGaeNFG7H8ilf0ycOmpO48hXOErBmNwBbxGF3RoW4ODYWwQJ/
UxiNix4RxdEUohNoG5TyNqXvXSnhpakOtvkeyTq2xdkWJ83/FUyLgEMVTGi6k/n8MHbrNMv5BSOb
yVJ+hVh5R4namOjvjJPUoPwnOgxI+sFAaYst2nIxG2OHTh/0aAoZfNfRcdzQU8ydQ2PCUfl5EYT+
Z3i9hW3Rjm1AbmiHlnbnmIwlzoleIkeWIcYwMrKbxUttcwkzYA3GqfeP0k1lDTUWmtFPQLJC32DC
WhV4ENKHDTjl9pp36GpqQd62ZenenpyYGFE9kADBXU7dBYKOHk0YOe+g1hwvGOb+hm/e8e3Ch/0I
FpSdtqV39M+L3jVgS78iFqgINQ8IAM34Q+St2FerGabzyYDFrxH/Hq2sVBDfhcL3dZ5THhR/CmD2
4mhgNATH934AQSExH/ZMuC6N32C0qBz+ZQVdSPDMJczu1V6zDe+jNBPLAJtUXmLnkl17SqGA0gPM
aOdQrWnhlIHujTTXdIQoCtsnhA3BgdWr3wo3x6PTkVjWoCaXwez2QE87RK8piR7lu1ryh/7aeCc8
qjHtrWQtXrjyZcYaWbS93iIxMLjiDCDbBsQeh4fa6SkaYPUqy8i33JnCwOmldBh0Ct5r838Z3/a9
iaKMsDRlxvBIytEKD0AbUBdh/HlaY8C3f1m1sMxocIVJau0Wgi1vpk7vQ5GrvrSxuGx8ELQ48mnB
GtcYDNgLxeAPEyj6w5ntn67nvw87/kwfkC9uGpMPfKJ11IcngBqxrhFVvZ7NOyRpfyBydwzV/jz2
AlgV0vuia+oIdz7cj44Un+Qy3qKtxCuc9+S0tp1ZG5pmW+VG9LulcBi7wuAm35XaS/ftTU8bLr2S
DtXrYFgSHDMIr0Xs2o5GMOt2HpsppHiHHx/uXFeBkdIAqeREcPY8vjftCs2oe5l7EeumA/YJx+YX
qjglCjLfggfUQ8Af6X/pNL71KS6aJYbzloLnjnkupN5JHZNOu2sy8utCQ7bWcNIrTYDNIOUbdJ5r
+08zVkLIyNrnJL/8Ycbl4/JpBK2HGsNJ5mJ0wkWkMOR1XXauFX558B+pNj3YhE79vK/s4Mh0ZsQN
c0b0prNrpB/0CC9EGx1V3tXqVCb9mqGChKC9jngDhkKoEsWlcF4wOdJXyQYYsiQk/kjblIWDE4J9
JhwbHid2zhzGEC9rRaSAQcm57PMWvl8+311ZYLHzEx0q8XNli5Q4cNbaRntATKk4cIzhgdedDIQn
dqAi616ffuxJhO0jC/aWK3wouiFZ4JtzmX7JWpRr6lDr30lY7WuJkrRHqVdhCgOJbUqaqmqf2fgK
fZPtyp0ePjshFop1q9Jd4pUlTTPLttjapjyS5DEfNujd8WVwmtLPODZeWmyHCoeMMVEtLJSuTBAD
Ded3sW9AQaJFLOrZ0BceL8Zh7pLyVvBsULiJSIkj5mOwdD+FfCYyda+69BazrXQlWW8ZfvCYomod
GiG8lHw/nmlxXy/a/8CN1xdHgdFwqHNoQMG1uSqfCxNyHIgWCjlVZ5dO2v3AXZWbdXr7ETafJ0Rm
gxeW7+L/meeUtTapSbnCtlXvJFsfAI8w3Nt3nw9w7ZBLt4dXn/p07ERArUkBoMKBygQ5nkUEikJU
woBy/1jG3wXGnEbZiJMsEyEflpQVuIqhGcGODVtlpFuR+vjvGrDvsLtDDnfaaOrL0pxkrOTu+Nke
UWRpV9CaFMBmISgMRZ5cYQ6b/X+AZnNUol7ZbefD+/cZjtnFYh3AMtZFUAA54LEYBhg2ppFTybjL
VWjLG7AzJICF4UCNL53AdSm2/gGhkdG0iAWZR8dnoiLvaiC5cPkuiV7YiN2MsX6hqiyUNO6E4YBW
G9rXQsovVmhnrllydMess7odk8b70FiEL867xgicy+CoKzOxFspi3VuhRIiZtv3nDYtWVn8ILA4D
brJGgSinaQTK4d/J0GoRgGtp7OVEDtQT2epnDwdlPJDHfNVXOj31Xw6lGwda/2yPDi86+yFiZe66
u0ORclHvUcy+U0xz4aaRGL63QwpS2AaGft+pet9hTg/fJiboG3EObzdmnXTKJafEwhMSwooozLzw
Bwh6FCyIplR5qvqLXY2YbyBgsANVhHmcatoLr7cR/72VdtEenHZhj0z0kv7wZ3Nv4c0UeIGu/J/C
MFNY4g84t89DRXhNWvSa1lg270jKWFhLcUiN6TsZ8RAr4GWdkiZZw/wbodvEje5vVYWSKFq8QXnE
+bbxTkDv7bMuPxSFWJ8H8BNhTfvMgbVI6Gcz+Y7AFrRYh2YnLetiWEwN6Yua1o5kDNgtj+vDfyUm
MO7Jic4K3q2grx8TQiF9Chd/vzPpfsMP/t0DAY5qSQ3nMLYeNOXWXwMqLS0B04pHx5h50TXX+h1h
iwOu4r/l0M3h4STUFLbZw2dHJLH+v+iMEI5cmjj2tajLCkA0LWqQrxw+VSio2cs+AkA8dUvMHLGV
2Bu+qCrNiccFXa0RMapAZOkGt1Mvuhh7wkVLQ6RR0aE+kP11hENbyWUtTJLEZuJfBRjNiStK5ZkR
srYcOLvRcAxOlikvQzdwRqfHbZzHROkZv9KRoph/saq9jBVtgT+wBRKUfWfxCPpNWo7ysuIlP3pp
W+j2zM4oGCcgClEfRPTHTegnPVvzVz/Nbasygt1SgH/WNhWNfnkB6pCz42tzW9wUzOBscVtV/r4H
VEDsXqgVGTo9aUqgKT8d9FtQ3QXYndMB2cW7T7tQdgNnI3OCF8683W0kPzZAnfAqA9Fl+OjAh6gr
F0sranvj2Qc7OBSpc4Oc5yg3zmozX4fkc0kDccJPsbErY51xAiOGV7XDqs33jHarTEkvG/43BxN/
yX9Lp3PBcT8roell1prMxhnp7yYoggrsvLFRGwEtambJzOKfzbrOO41JPFYuYK5s4tQzxZ0xkNmv
nezJWU4UPHqo92K+kxJVRb13N+rtkvQDZnN6s2ADro9xA5XGXtGboYgm+YZrisltxYS2eHJLtM79
8gSA9mDOsGvCxgS3wX63jtKFTFUYTilNQXRpkY/RY8rwKmnubNbwIdc9CbhTyRJTOJzwUrGwbl60
bBJWnYMVsZ+NZfIpTaNMWASNjG63rBFu3fN0ZurXaW4hshYlBPbQz++i8tXQd4j+wj7hH1O/559f
LWswAYYKelaKr17l5RvwN9psWXaSGYn5eO7uc8SuSmgmCuyVttaSELI9x++enpdwVgsWZaGTre//
ah6rqmurCIbQy/WTaPOOX7/bKCQDnlNon50/Fn3lOICPGVkyKSYa8qbJO0ZoLVOTBoqyAzgTqmWI
ZElPWAR0hIlxA1Xni3gf9hULMpVMP/6MV63NxLQRTQR/34h/sA9TMg5UOiuHL/16N0QueQkXAhkX
kXpkZw==
`protect end_protected
