-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AEj0Mvpj04XRw5Qp8tQP/A1uHL2P1cmAG9RpPs2WCGM5BCd5U0z7nKPgCpXo3qazMD3mutOforSZ
kjnvIjsghwcqkRuCfmpCztaKM3UQq84YKnf2a5su+eybc50q+jy5GbdudzK8EhWUKuXSLLtwWZOE
3rzq8+YxMH0OULksN85kImhBNv4jOrgA1RrlzCtKFPVddpqPQiAPXagzlsRzlw7hECbE7+eszrw8
s/bVK373j8AemPhR5J1xlPk+C88ZRpTFriHKYAhC7pg6K/RjKQY3StxBgAhdK1cfCLehA7z3aFjx
V2UTRpD2VzgTRMIXule+i9UB9kM3u83Of14EMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11856)
`protect data_block
RVvNTC8347tRll1UOXmTmMUWZOOrx21E+SpwNIy3Ypiagriao8euCyH3+BY3Y8iDSOScAhIroF//
TYGrEdiKhotHLPxnj4a398hD4SXPRz7M2pM0h+u+cWYj0bV2JgZ/kqBIluoFy1UcNcU5qSQItpQw
nGkBHKQ29iaZXo+EBmV/EpIWNgOBAq4k5EY3qJHRR0IIoD3YOaj8inoUQT94y3ho3eBYbpwiXfS/
3BHtmhU83kVr94CVWlX/iel4E+yYomB14JUx17l+ycxSpmBBSF03fl1rDk9VPEHxxkspUtF5zU1j
tE8P5dm9bcBjB50bbnnzWg1+Q/TVB/sEThA90/pvqIx8dFBorl9oP2NjTF9clA3VmGyKrVpDmil+
PQjrqZ/aTlBOvd6xuVoYTo5I8pZ3xUdTianiMLkf7yCaDpgRAXdIS0HpASmAbRTctlpzQM416pY2
xxv0YDt2BTD41ZudpVgqp2ILFkVX7uAJE89S8SaL7sJ/l6zyDZi4qxNJsxutilzlysZmPDqRWJ7d
6a54fSLyPW4AVpbWTTVCTCew7AXyGcgNTLAYoMY8k6lLFA6e9QEwA/9p2nKZ4jTmdpJF6fmMlxx6
skBLopckpSZWZDzDGdrrIU4faQqagdw4iOp7oBR5uG9Vrf0YyfgjjxG6+jQZQ3xSeNaYnjzrxYyq
38VV4O6t4MRz/HuOo4lqe8uVIwdkgaQ4B/dPv3Lya9DHRS6AQOTrjwm8UQ7baOU3yNSWlsRkpNag
A6L2gQf6p7OdlXwevWxy+wpCGtJsxq7/lyiAsNkHggDqm9nnUL2TysMFhivWuv1uOSMNN0L3qm2u
7RwdyrPbN+TsYMtnQY6rRWiEORctljf7twrg/IKTqbcok3ILjDq4JxTBw2HtHWcf8X8R3LTpjaUo
KHvkW2Ns0+3WWPTQ4SnnVAXHFonqbJr1dLshIy2EQ3i42DajwQUSjvCCcMSClOjDj4TP3qSx05vj
ZYdm3AjW+8z+tAmmX8eFtjp3S9wdASA1Wgpr/DdQV5DsrZ58lQcp9DLXPC2lwOiGjeUn7FvJIKGI
JU88eu1Hw4R2MqXNQ17VmXlHH/a70e4/4LLt5OA4PDGgrMmup//ZoScD58j9jrzse9FN51B9yA8c
qpzFog3f0cnT+ja6qgaoe1W9QiDIJ6FeAC09SU3m3AmfidtF3AaIOrnTN3GbSuNtVKUX8/Yo9lFO
ugK+IgZnM1ZOFWLl//NPIkx7Ba7dAn+nzTtsK0vnu5iLH9xc4pkHb5060eXVrxdzqducg6PKwMnO
KwR7/ztEKjv5UGdFctcOvSTKg+89KhKKTf1QdNxi7bILw1PlmZViFapWQdgG6o2v9nu9EEkWcqA5
AMqBOB7g967dFBebxEeYmkaQKUvj2fW3IcM1tVYutsomhOvetY8k8X4mGVNf//YCaR8VGRPEeUjH
vyX7wrlwi8qUfJwa43TEzkMv56e7iBAZg8To5V3ILnBrquJmf/np8DaloGOI+ONn62/e4OuEaLgS
GMlSEEqxlFuQZUz7UiTxAXy7Od64/eUOdC0mfg/FKSpLhUjZxIRbcorIkAZHq3Us9/7yIzvgOgwH
h9O+b4t+V8a9dmP6r+rjHrLW2cd6Ap01kkYzEdBfAxq5BEpWl3ta7L6W+dP7nKmO75qSyGESrlqE
P7gT9i13titk406Yvuc0Lwf3CEFK2OAOSCvUk0iJUSfKltHMeTGEm+0sR8TkJko2lUlweOX+uUat
QAKd1ewknOaBlJ6UkGXN5YDZSX685bxyr/Btww8HG5rmmXYjn78di3omwNmLpz48+U+3QymaF4Xk
q1IY2T3b+92lkE+Q9vvJ4SUPwkHcGd1htOv8rLGM0ULemxU3vlO47Jf1G9LG7zs5PTYC8I3FoSxq
0tMmCDTV3hk9sgec4ugP8n36bMsXW94bM1PYrPmLtMZLyr2T/owSVIVmktw4jRO37GIE4K1QeZhW
Ruc6/Av/GF3/uaRxS7ONS06PY2FgIoXuW72spnftNaYuOGYfi6lLONZalRegfjT73v8AZHuW6+aB
GRkkz19zxRs6qA2jynFwDNzzUK1YK5xenSUNt1CXyfBhlZuoDpyQH5oxZnXoB1bP48LfYDFUo3Zs
wC9TQTTf+2DYSsZQxQacp4Q5J/Yev8EXvmhG8BvokQoIuHXRLYw1KPHc9zsePkAtS/1O9xMXzYTG
i+8ravrjilWy/uOuC73h2p1P3zT/RmEq/nqVAULcFMES87uGk/EyBvZU/nYzPP2JTJ5xtTRpmoKz
J19cURyG0gNsVE1AQ56Bhyr01CQYXD/buLVSS2LswNv3Ok37iz/XGgJ70TVvs1oZoqwvXFKH5PQE
9+jFmp3ZBs9ZyBl3ZjayqakIivmul2CB7c+dA2wFkoX3JRUpzOLDT6rAGcoa3J/d5AQ5DHjn4Gri
KwhDcaNzRo2CreQz+vvyacU1W2vfC5xFBCcgJkX3AatJq+fwfEwzYw06qEbjHHBZNc0EMynP+z53
LZ4MPfmQYgrHHT4lsvnbBBoYGzxX7qL5FLE0yXJYyNxaHhsCJ34+UWaa81LpPHA6pTTPbpsDjMJw
tVOpIbMuOws4WNess0sCf0E/2WtmN+oAVqyaY4v+ALHHhffWazev+SJ/I0rYgpdiUftdCJjmco28
ptx1w/sKs9llvprZZqkFKDaynTxNx9U8j2Q6det+uymIMhGbCW8Xv7jYwUb5GlDe6z444MeCW5yy
hQWxuzUUVn+ZBYLsWOGvXPa1sZ8dmj6PkAhoo2OtmO3/X96XrCF0i6fcPTGDi98VeDpXlGQpJyYu
Va0m9Xiv9MbrqqY1pt1mbqckWrj8H8kLulVAEbHDA2r6flq1YnWpjw6J9BYhba/FZWQaPREgjof4
Y9B6heVYwgKr3RZOaXq8UoS1ST+C6oL7Dgk3Y8UeaI21ai69yxNJT4c5kyZoKeCfQyinw4Tt6baD
NPe982G3COvkbxHICdE16Qsi0RdUvjh0YmFhUlKQqobCdzwHarop1ut3tfAAoyKeWN77TOYs5cjI
MGXBDDfDH30mOiUR5BbdsJVCdkTWQkwB24MrMKf87g6+xlLJ1Sa4cynBIXZqpEnSD+l1Ayz7jDOp
Hq87AShSVmL1b+rPdSBpU3tKiMFseD3ZGlkdnRDuQHTnoflQpzumjFn+NGoZtOB8yFSM8mvgJMh7
RWPhkb/JjVBtU7Rb0oE0XapFs0d9TRqRu2gA/PtvtOrtQzLe54RQuedu0tR8IDPBfRHZBHrnhzmc
9cbh5P51Jtq2FPFuc7oHjKDRayF2xrrovuQSZ5t5Z2Evewn0aX+S7xX7/OJ33d+zk7tWyjqquqYy
OxPU3e1JVGvpb+LX4waMXD3qufQl56MrTqs6GHMDtpuHeoT+zdn0WH7IUOVNkk+by9ya+R4SsOcK
zcmRgNRf0IFOyfB9an4yjprf7PSGfETf4qP9XydExYVNqZ1aw4e5KdThdMMzaddKb9bQrmFG5Dqp
tpPet6fFDUi+8T3J60IXA6qewoXFskMGzSLphWdb0Dv3MZ66PGXZP+hhcC1pVnW8ywoE3BUdeNyd
7oczyajY0lcMTStGtT/oUCnzWXDpe6n5WzhdSW2rCGF4WqLNHEkvjknvWjyT2521jsvlFOIgF3Ky
+xFbQvC/CO/StLe9Su0vyi7kT9cH7j0EkEEJVNkqTNGMuUDYfgxKNnquska0LsM0SAdPCrzcqJZ2
3FA9a0xCsxEspA14dYaaoCWBtfb3ivUfnolOBqk9zIVXprRmaillMFJIVzKQngR3ROfU/xfF/i76
9dobP4dboIOHg0iLqmJzcDXeiSSAdf8OoclKvF8ZrvRLRYeT+7NSyOhR9ydoNorTS17Lu5PgsCOc
rHwE5DsJnDfsgiEm6J5bAmVzKunpdb5S3GNVWs4V+EJKT7hH6E6wSyaHcl6z8NVdLlGFEofUhO9t
oeje4p6yYWP9FO6MuY6U0OUe82oGrhnl+yy8a2VAgBWOCxiRbRMs1kcoBBpw4so2Oj556YPOo7xc
IfDPZGH3YVj9qFaRG6vkQHuAPHfKosS0QFTr328Ik7YU97T9p1VyDwzo0A0mFtdGzZezD5n/rChG
cSkpDR08NynCVuxFq0vQ6gtQjhypOBjWOx5aP1esEhRPZPe1RtOTC3CQ3HeIjbqNpHy/dRhMiqlx
/qYSqksrUkiMdGuypDPZOVfyDksIuJ5azoeLycjjvXXZ6Khiyxx87Rq6D8Y6hFFgh87ZxBXqtqwL
rjbt5bg1R8ZSl3bDJf91guIuKryYuOD2yqZwjJaL54RO+2lS0fRqpltp8ypnYcPG96cj5ZprLYrV
5XtBiA2NGYeXAp1ulJyDWxJIjvhjIIOyzaAYG+suguiJ2fnx9aTJcqhnIEvvWUT1q0jyOoRYVmjg
SYwFn1TYTUGWgYeGW9Yaicen2SqSR3wGlZ+zXCrjc6lO3l3hBHE7YIcJzC9abyzQ4Y4DCaUzv+ox
g/ESTeTGZL6zZuGrzq5eNt6C7uQeuDx2IGBlAnQKWdC1Z3WqiCV3vXgqGfOdLRNKArQteBXLKmGk
ITalsIWEKkirbHoeLWE3+MhGt3vcmxFAvhMysZ8eAfCzzWb6eUyorP6LsvtdGHQ5Qum4XOzLfIC4
5Pv5K2NLaBPSIzIrZlr916OmmLZ4MfZ/P5GRQg+wYRHhqL42Cqmne0GdN/3RHVE+N5gXdoVIh0U0
usOdVJhwn1H1bbUUDJHNfimDzA/AgJGTaePoNvKwnLFdr4zbKJNtOrnYLbwQaJ15W0tNXVGO92Zs
yUWHXWhi4xUuIMWCBOYSt+X7rV+LwAo2dH3eLwnpqab/I+/D9ClWoCvEYvbBW+0h2scSChDoyyf2
y8gt2YjYNTUo4aMlXgQxSr+Xv04c1CRk8+rweAkKySj/b/bJBClqMCT5z/KHKAibXeABD1ga5hUX
321jk+XQasGpfUCpvOi8Au6eCoXd/dK32oykQBbIaadrKSqpqV2SGNiGs1YbVc6iFGUFsgmdmWbT
5LzyK07NvAfKhI3HQaeKZ6IokhMzjkcNC1nnxchqICe6lhp3k4bny/p7P2NEP2QYHgyTw5OzKPej
XJ7MQUoooitOfz9fzVbhHW+f7aGCjr9XIcOo1rKu6gdoN8r41CVk8fpG0/TNcbwS+T4HQngQienz
0X5m7oTPVbft/DhrIS77W4X2W5zwKG4f8cClUW7C1c+N7cIvX7xeNzK6RXNRilQm7EaglF+mE6GW
SXyiMb5c6I9tyPKKK96T4ZjK07JtHA/yu52t3dTa83AIRuNK5II3rs5RMcZ1xokIbtgP9zwjuQRP
PChXi6EuGF0z/pioafWxRRj67lRmeCuvoIEUgD7+t45tMkllr2E7uclVdDoW16yPDF0nuZUoUlT6
qFi/DHf4xaIU5rohnvXcQSkGogG9pPxjou/Pygj0QXNWtMYvYWw6L+CrrSD1yOhFUQ3Iw6c7Hq68
1FPN/twwjjB8VJ5kDSmG516n8Bf9sSihzigCxYXNiEYmiTdf7ZshtFMudUFcPm0KD5s9NGQ9DZZ7
FSY8GZypj/j7EmjvCm1dcZvwJnwfl2GGHeU8Fvx51PfNXCHo0ZlMMVJnYcqfLv+uZodn0A6c9zgL
PSCxZJs3WJocKZHM9ZKmZtzrgSQE7FgQc/D7x+4+A3cn0oQ1IzKXsn+8nKuj/4g2nTn6rpaB2csA
kOI4w1/PB3AMI5yVf+yjXoKlz1k9SHWiYnb+FV2btYyGT9PA+mj54auYdSP9hc9jKjcg9q9YuGcT
B8fdC/GVe79N85wZhLY095GXv/G0ZvBoPRJZ+lssHK7kZip48rlCUAoerv6VGWoRogTj7h3kxUl0
V7oqDxGw1VB2lZ2uzQeEIuxAsyqdVKX/s8yui/o39GeiDlKYeXEEnuyKQBWdAGFxsFg4RwiZfuBc
foZP6H2RJjfeOSxqZzpmlROeL0NXl73SylJGiOE9bdA32HixKj2vKqX/64AVYzmnYPguRtVZTqs8
0FwX3X3NZOUPk2kCQAP7umt24Nv4HyV9SbZDBOsX1Dhv9uRfNuXTTDzo7ePP6TqIeh3X50OHIqtt
UoXDpXZKfmcuMUcgb8LkxRmwYpHfMycA+YurywOUZnfN0OMkwoQVF5Pg1Au/fJin2t2C+SJA85rC
TNqHxF5BLuaZxpOmpQoiQJi9OhmP/wmN6BjjJfOTLQShM4mo/LGZsnL2EwQ7vDVxKau2+bSu+BI9
YgzHdUu/9aG4GlGyC07Yrz5K8LnKWFkfkMkO3CIQtKlUsVuQVU7HVY6HxWXl6/UpCnl8PlaFuOnb
Wp0kNNtChI7gZhRKjWWKmvRIiquLX+EjsvqZFQkqfqHwk96wZLHWKDhKjocQ05wsplsVah6WsOZ8
gUkwvN2CRjS986PjnLiIw4RLXpHoPUFvJh3DcvG7AurEmv4UXn7er7z11JUfW/7ld9xDb26ReisV
Rhsxb3OeSyMw08em2bgIX01nQTkzffEUBqI7qkORBJcP5NFnqpShoNoeKkTDGMO9IY+gM6kr8lQX
jJSDbo0nLVX3xJ1GC/i3tDj5T4JPloNreQ66yAbG0Y/2rotetODua4rjG4Y4s5XkNSMemQFKj/l1
9BASzs9Uo4f/vHwPqgtZiclT/38Dv/v4oMRDHkPFo54L6y55Uu/+b/SUTR0bVusr/QYHPTj7zDV/
ezhwmuAc2kcyKtZnDk0wQ29ZFi1sqqQmohmJ5lPnl7ymT9aRevfxRV9y6Sd4qvNHdw9QgRPPuCvq
+MkC2Et5DUOBfFHjYR0bgfBRvYHGIJQACdykz3FAtXf5RxPlOrEsV8JpSh++SjPRZKdD+fl6ZieC
8DiJWML1k4Rx2Q7hRjLWX6n4fe8XsHNyroVtdbGzBnmL/RJw23K88vFpEFJkqYYrQLtgAja2Xl/h
p6IL0U4idCZ5aqXX98BAG7BvxceX72KI3mmU+qT7tfNg+TpZ7n2KA5wL91B63aVZDouDLyRcxFm2
X99Evgt1UNp5NjprfHuRk6TwdWq6ow/zDdbqEaPsg5hpCJPB4v9Mda2u6x7Wu1p+rEnlPXoHN3ao
Bdu2kCi/IN3iZya1n1ErrbPlaGJcLWaG0CzR7U/qSF16Efo0krhTpWPQzN1P2SDV4XrkNk59klpT
PhUBcmo+BAP7/+kkgrT9gL+D+IbBvpOKIRlDr1mCS762UC1kY1CHF1AanS808rL6LqWW3anlef4m
1LT1W2jyHFhYsAYd5k0DOxXYrPyRY3/IUt+YLW3VXy+0dA4JfhJgoQH34EZ4OMeOGCIDFOUkFwA/
vQUGgpS4ojv4KGieaeY8OJJ1UnRJP5z0rXzHTBarlvNIlKnyY8c3o8yp1ec418HNCrPFs7RHQHNy
4/Unsf1GR6Am1imn2m5fbehh1XtMt92kb3ihy0Q+NI6bkg2Yy8tOWIVgNroPvKdt0aCeNB3A1klA
Lsq8YXmHPmPB3QQCItEJovunXZdZz96jA8sk/akkiJXtSaWjHQT/gDdvIyCnz6Gv10NqoGSG5p8x
S2+qZ7GizCh2rtNs5dl0+/sewT4azt1Wy3JloMZikbasEcBXUMDPtM0BYXCMMcL5HwCfyixHmeR/
x+oQ8Mwc8oZx7p289WUMJvPRb1ipt2uZVR7t6XzUIDEf+KKo3IdpZPs5JlScnIyBdAR9+RwkQzy+
srF6QwNH7p468IrRCuMRSiDUglynrgsfwky2tshX7DnffOWim6YS0KV2cNvohf06R1E9ZoEaUK/b
Iy5iSq6rysFSYKVpllJhC5IZCwfLNfUtMF6JS+wswFJz86polOoItqteAs2y0yqgiuXTkDzeYWUU
JD1p+bQFyjpcBMx9t3+ojh4h2XqtNTYH0LBrUtIs2uZjjHHq7QbAtp2x+pt2EcR1fDIVGO2/dGZc
KSPvD14GTMx10I2J1sydx5k2NyCHhAwq5gf0AkbtRTbjXkR+GoaiPsCf+OpfQHMGRV71UjzF6lyu
gVptiTjh0mFrq1FI+Go9cCGq8l2TlvdDnmrArQQXotTDIMnHDypS+iB2R1f+fgoV54WJyVUFweq3
he6CQdw8f3SNk+SuiIV2CdCSzHbMt6anAZBuM0Dwa30X/XNgduIYxWeyABVsA8a85Ew3irF+pSsb
ATFNhjQdgTtPcQ7Qd6lqZUlQ2/v/0apW/dNyDm99ZONTGPGnc6+KYU+bqHU+OkE6vOrfvfxnqEE+
ZHwL4FxM4gDzHDI8XD8ZGtTAUXvBd1bWpwZ1BQG/MeLxDBYlNR1pD+IByuL8IVpqSysXWIKZAGI8
lqhky04FyhIvMkDYJK0YVsUzmq8i6smcJra0V/hUha+2f2uYCAtQsDxQ4eJ34JJ5knl2qPFUtDLI
UgqZjMMbsp2a6+5DXrC60a+NNIH3xRv9cMfNTWpTFkaLE+h8PLdnaJpXJJNWBKvvMpMLZjSNGRWX
jbUD3guJL6EzGXl7kQSyQyj+CIsenbBegwxSG+wnpmpzsGjTt/IW1uqPk6tat3WQcZxPo7pVWyZl
8f5PrGXbrLzwz7NLUqtg7Jqc2eeciKxD6m0s5mLz6IM3KVP6sAn40KCaqGvYOP2ePfYGBTWxDZDx
klNJhiRONnbCpdtywWKgurFPOH1+9zopoPBDE2l1bMxQMJgjCk48o4cmEVLfRCFGS58HbBV4Pmh3
CueGmQoUJYhwpBrBvGOBUMdIWrTTziw457PHfr9Rz6M7JPMUtbJ2GJud+f4NTLExRwol0ER5BQKI
V002YhDyzTSSVsg/Ev4vtLRCgIzsv6d0YLzGtdP/A0gmx0na7tXFkbOHElmNE5ES2wFCIrR7rdbB
D4SW7Y7C4l090bA/SMLvqjhTnwgnTscyQdYnYIKy/wIg5LomnfaI5KqxlbREC4Uai0/uW+7nd5eJ
K8uweYXSkbFgWHlQ+X7yIwOWuav5ZfJAa/C9OxEwdCh5N6xNNbHui7eJ8V9n4JwbShh2/HTjlhT0
l2PPQvjGr2lHOc79Pt/BvD85QeH4vIOCaXT9AXgnVSME9nGibEpR6YXe4yycYR/KYvktOFXv/HUB
6wFCF+NZnOf342ZxDtuT633hwko0sIK7+Tw/r8etdI+NEPOgqh3qb0A6sAYJylhK5KJEVNxDYqac
Cshv7KjQ/uzJ2K1wzxiIoja6m0b3SKeOl+SLeyJpomrJU2gm708ZO5yG80Z785b0tSvt8JvhcNKU
S66yV/mSnDf8fNdBEudnie3tdBk8yv8elLgiYFJuK8fK3ZmpDCZD0kZ/Z5haooWhPKD4B6pDcB2s
zqcovTRG1iWQsoM+xSSoDpALv1P4x8NA5UvNyHshpVFNBXPR2ZqJpaXDtJ2jlDP1aGObJOBDQ92c
/+iQRegVSMm+KeLhgep6BhaMH+QGpMCyh8/BkV2CVD6c9SA/cD91TkqhgW09Vs5Hix8otzGocwUU
mMATUgDFF3aDbMHpAu1wYuSrYL6o2PKN2x1fITjfsFAXLDgy+C2TNVBLn0vJQSXcP66ufZ3pErxC
ztqraAK0pns8pRvMVliYCXUpBxTdGI3euULJF484z9IkQC8At/MueBwF5/WuhDSIGCG8INoJYc3K
RUxvh7I09augKy90f0fL8gRQg4mWEqLGQSFiZ3JHPcW0RJiGBw153vXYTjkmO7/dlUcbzgmCag3g
spaYnKOTzUK5h6DKPmyRCAz2+XudzI+mDcKbQlIPxxHV5dx6o9PXSRH+td89OF9yguS/DEAa5z+Z
zvq1vy+vigyl++iqywYRT1wDjKQ0ULpxqd744l+rWFoYGpwBo10qj5ea8wkVyxj+Z+mEjOKAZFwl
4md9qZkLwM9gCzvPBwsYCfMoe4jLSvpkB30WWUE55v8R3Snfv6PiayzopDxpIHl/O9krmSIVCY7P
QsTmEuRbg4qnvJmyOVh2XX20jXN2Tdp7IRZnmYRomOehU1Eoj4C8PerXLR0eheWgS2mJT+UolrBo
ywsgSnDUD/PyqPT2Du1jqZcMkWEzd2PgXrKiSvgQrpPClBDMIRi8BXGNadBMcVEIP6fvTrEa/lMo
bixGbD7GaZAZ4DTnlNlmJromxHRQS7kS1lj9BHhIWtRwNDghS8vZEWZGDeFVh6zhfknXWhA+yJUC
L9ykm0qrQvvfQpUYHUavDWY0UVOpsdN0SkX79BAoftV5rKAiTMFqIulLHECvk89YGX6hQKn0rpCJ
gf2SWKmtElOuAOADZ1VGUGrbAdCxBTLRydEEU/c6J6UwykgT3vb9kBAqcMj4zATo4KhpPKiQ0aDr
OT9KmggkjRzT22x+JaYTuZBBNarFoij2xMG6JS/H8ytci8SfXN+tKotpnLAatsOPBMA9ONJvoJs7
XTVFIgJvzFRiv08qo6Sf6f39c62OeKvPGzHHwIqX+624yH/5BcGsz9Ms2HUirMeJvPtGCZGgA9Yd
P/TqA3huTMkeyTvnHYnZwutj9P45rz4yRryYahzN38StjMBEZ7ovOZfEFi+hj3iyRS7LSSi5LYDz
22oKvLeTLSrUi/lk98X+F2gOscUvSohrcswXhLyc9gcKN4czqNGA+DVcKzVGxl2wDUuqir/EItVN
4TKWE4Ya8vfREqDPc1mjhoe3nIFDkCceQ9Bio6swJcAWX7e4SqtI8rfK8PMKZU33L6Q24ZE0gjLI
Y1POo52rApW+Ss9MJFLwZu5gSgcqtwksvO9vClwqG6/DB7s1bxPDKXMp5sjiMpfIyPmIvhgFOsr5
RhTieqKvNBzP64pW9NMYZvyBvhyuOnIpSnvilJacQFj+U9uS1/sGNdchYXzNfXgqA+R3H2TMBCNW
fv05pGH3CYpG3cwpxTqwabRVQAfw6T+QM66A7x5UHEP4edGSb8aSlw2C6s3qqMJbJNGOVXzXXMs1
NIFs6fU/sZfwST8SoFEigjA9B0/sRqM2A0AeSHEzGQNuhvCvOkDtYUryfWeRL5Ys+IY98uir1+lg
LFfCdRiT6z5d8YFScV1J8ar38hSk39v3Fkv+phH6w6NSc5i4nhuTmMGCbZMKSyLWM4Kbpcq368tv
NCb75b+wV59k7FJx8I76OIyawWNAZdRqY3rDNuzkzBj+F+Ik3Yuc/pOv0wQRXuCAbYwsiGJAMCbv
9Ut0TW24oQ39g4s1+NpMChkCd42uu6CpUUXt2VChe+gzw0OSlvDexNlq7PlyGdzDoFwvLezzMADZ
rFeXfI/SdIMRtRV/Ujd53KPwl/FPl1xWw2W8ezm732xKP5HCFuOwz8iZw1VDUJqrPpQqekdA/6qH
R7OpIgFn+5XqjBtDr63YEb9ayTJZ3HMBf5s5p0NFh6eyh30fcYEsr3eAlUsBhIORrEAbERx7J5ea
+OQ0XvlGxJEWDtk583IETNvvyJXOGyHjop1essCPm63ljmJE8W67dbAaMhbMJNc3aAhwz9MxA6yF
c7RCW34CQz99O4IEYxyeZxuqDmA1+lIV1h3EZtuH4A5gXXvA0nuwJn+1d9pRb0FjOb022pc1oZ4k
znX2MT0PgSSMeyT47fyh4OyLy7UnTju+jIlB8t+gBW3FxOniMGIs3SVQqluMqleyomR4MYNPIkCp
iMsfgDooiFEo5KKVzRCikvIe8zkMUhEFd/wHIG8aS0CTKLjtHgHkuAuLur/s1G9XaQjMFo7EHR1O
Mz37FEwYtVKKyJItr4FRLE03YpGePxNev9qfUhr8NiqbzZ1oelJq2UgFWucRzEv5bVf9Hhdnh/CF
92lrIuECE/f3xro4bEHDZyP+lUo8rhnp/AosEmKHtfJnLkX53Oc/wfUFR27ja8D5Vq40umQc7qRJ
hXpB6Io1JS5FrkxcvZMwWSBFddvTLm5IS25+jaX+umMfUD3opcyFGmS80AwbVOd2rs+2g4BmDZmu
KB86RA5r21nGLbLf3UkVpR3NR9rnccLBg4sDSjj0wfoqTRBEAP6/NNADB9XBJOfegZ9txaYgRyJl
zWOvEvwo6j62HdTNpXT4GKVqGz8jOgA4xMD/Z91vFmBsotPYjQTas9yDzrgzPdFvb3wUuLU4sGuq
j1WoCJB40uF2Yz8x9WYWPBuigSmiol+kx0157oQMV2BM1HZG1lnsQPBWNZm/zLe55SIaQgi6nUiB
CDA3XZfn348hbRdrrvBMUSlOOGNrNlUz3NzRfVuS4U98c6tmkdulw4ShRgvywHvPZj1bXBiZzAuK
BY3lTUU89016kDAQVqhdW7RH0R9GmWC43rr3aL/yqX1H/7uPb/AhL4t421GuRPGw0Chl6XDoBx4h
CHnZ1r9QX67L+hfNrpMIPvV8efxy6vQc9kUklZn85+kz5Z4vheA4XTigQSfK/vj5/7I6C6buM9PY
NX3TqdOpfbIqqjqJoAVSJ8pt5GXxxdwx6Eb5wbI8LSN0Zzngx7pi79HI5ht7ZnUZ46ouSfMCdYoU
LvLa2OzKUEu6tNAtUf4LUEtcI+TaS1QcyeOwSqc6lAxareJKgYbgc9vRmitaOGS/8yYKi0JimcHM
fTlLL5AGp3/TXLTTBye48vFT6vanVhUKAYIgvHjmjjxbAKk6VH4EImfz1Vv6q/c3Xfuc9PehbEFZ
YfJGLRDGyTgH6wkxyea5VqJ/jzC3hst8J2UClRPzKy/Jsv2K1m42AsBfiC/W/YZ2xK8JHstTgM9h
yVc7G8j4wdpVa6G8R5aBdDjlDOHuGnGVO/kMW7bMcIAkwGY1dDax08X6XXQnUQVML9f85+C1QNzQ
KiutVCBW3oSIZn0xuN8CiDtasaBalPENUJhe4POTAPX/Yu9mJLe7wwCEHY0zafEAR4HSXJCJt+x6
mSLRjC/g5ZRhUFDBoauOK6PvBSJPt88gFpipSu7AFI31QHUrzGc7S8wqbd3+FW+8hPPptW+Ia7U7
ceVT9wVJBB1M46ZgE2O2yqznI6dC8k9lUTxdYnwjwLx/rcuO+9KMH1MZk7M6Xyk5S2ZEo/vQW/D3
26byeDCC9YAK92JZeA+Buzm1ty9dwAX6BPsnjwd9mHIdzshIs7TnnH4Kb0NVN8LLdvfDzFle3PUs
R4nqT1Bpm5G3MizHwyywMZDM123tv7Dx+kJMaXuDHZUyb0nR37FC4uglxVzJHOzw/egPn445AA5o
FR7rvlsqigHGhFjpnLgYrRt35Vk2G3Th1IHcLG1WA7NdPfCgytD9+umdjRYEwVb9mGnaWTa5icgt
kf8f8J0/FqIRi4JeDSyItNCJHu3xO0H9sdlsF/U7+FA7H3W/xD/dgXr1CJ3DTBS/aWKSBBYJIDz0
P5WHxDde1MwTsR06u9Q//RjFy/nGaVJSIjdhNKbtsXQMHlkp4IXyEBG4UX4r2kP5yQSq+l1E/R34
Swof5/Pklq85ULwtdStCb5tO5aqr67uVSbrITThlrFO2QGtGcIwVcCBRs1oH2ZPYKCEP/yBwweIS
nStyNd+rePhNVYBjR7onv0QIBksEEv5fKZ45zBeYLhDjSf/Qz59cXemiVmm8IFv56IYAm9uEY7h3
eOqWuZ7TRDkFXA7AVtrAiFJUjJU7ryhNRYFMc+FfXU+2Sb64kz8bLm3sK+J2Br/RhaP+C6lMsj9e
zJVWzU8UgW6iBZ3nfcwyK61jVwL08f+Akumsc3jimjcy+0YPjhBKZc5WzEn+KN1zBGIwaBZE43Bi
+I6RDwQdKA6XjtoWdywqK/ZC1sartQTUNs+zVhidKMuwyR6z6V2MzwJFd54PQm2wzMyXCaoEJPlg
mdtPMK9VJuifh8IUK9SoauAZGqD/KytpA+cs2YjhNScbAwwVGidrLECSMo5i+zZsDqTUdtkyMEPR
4ql1eF9LWgGdHrgMcc0b+dCWeIloxuVnrc06J0g56kKYm7wOIgDna1HPVqNmLUhjcEk1sgZqwExL
93n10VSY8rVi1ydtaCeGx9jZMTUBj9LXkWsjXy62xCv0lKDIr5ZSzWAWU/G/9MJ6Z39slcdHttOs
dzxYLp/GQWq1q5JooXgSi/85HGGckxbaCjfOjt3eulIeXzPhAdajCvECvOyDxnMJNO3oRN7gofWu
GNQwHdUGGHldt2s8IYbYF8DKPaYfG8LU9Vwntidl9X96sv8XgIkUcYsvN5tGG1Z1VPZ/NoHKZTS7
JUiwCPtqZ4tnIelzOmILamOc+VN3eT0EV9cx8Fnb4szGO+1qL4hwmTWN27E8CXgfGCRlQyKpaxxW
1RTFlg/3UIj4cRoCsrpN74S4p5HMFe3DtxQEBIp5mbJxoxKrxHZrSbuki0jlpkU9Su5TF/0Pe4CT
T3+Tn5aM4fB0PGb/dv3ZpiN45VJpp1oj4Y21HsEPbvckLnAJ1r+iuEvbTrNQRuZ4whVN5WD/DOor
91lcsDbFBTHvCAfbreigyGTWK8B6DjW3pUhSGH2o2YdgKN5v7ug7CfYq4ejLICeFbwdoTKqHSLRV
0TX8HT2mFKK3kXax9++DrD1yFtjgMYTvydQhzQycam5lIKlH5shhie841KqZCK7Msh5OZD7ftL12
oW7MeYMinHmaj4+KbjPAGF8Qb3svGqnruInkOTIx7CUXdq7/umucCGGQftJpMKp924An6XJ5ZUQM
U45HvxNjl8Iz+khyimOslX1zQ3A4clUoQ3KRkT4rHQT3Ygpvw843wLtmuYfH191uM2ceqH/zaelZ
zBAFO+VrqdC4CCahTyJ1NuqhURdkyc8hCRYIbLgQAeRkkvEylWTse+ZJRxodprRTq3shbScyvo1v
iG86cDlXF8PWKfMBOl0dI9FiTbdT6t29c7eqpcHwWxX30EpF1b1Q7zjhVuOYsoaqQeldtXlxr5Wh
n+nOPxCXHa1cMwU9QvLv1DzusjFRSj/Gqe1BXYJFwfH9xe4cOxqiTTmcrEGX3A0SYDgDml4NmTSD
rFX+9VCm816LmzmnpNMaf+o62KkekJJFBhk6FR6wCYt9p8EFf/kkwPL7mxQTZp7l9ZnywAgy5UvI
PbyEOId9ODglA/hERY+jzQCUM3vWpf0IBENNFqEsadSqIyj5lvITwdxroPKiXt5le109A4vOPYJq
jmy9lyX5TcwoNUg7KLHCRMWSVWSBlNKv5X5LIBBbaWCWo6eqqxdBC5/cQQGH7l4tz3WVGeCZU4Vw
AxQEPbwzZK+rqIpnRbTJEPdU9fHmP48/RQb/l8lxYroMLFUiBuCkHms+S7MQFWG90a9KYS64Kln0
Iw5cauLK6dIfiPKOfGm8t+QjvWSHvAJm1E8WIPXy5ST2eOe0htEtvIawGUYLtU8qv3NcmOupKM9f
Z21A3MNh6/hCNM7hnJdYG3+8mk2wJxWGnuK5y8JSNupcg8+k0CPwBG72/urtUpd/y9xCQpVjeiKp
WljOGs00vw/eThNNflNJEp1JmK6oZfuolxDqbaS2ZKGZ/dwB8U62P0LPmSolt6P+pETmBdVqnSzA
QT2hIn+LjS+LF7Tae0L6ZxxQzGkSoYnpG3h9C/MGXArv9IDeyPDfUptRX55gtEl/U1+LcTZnoL4g
Nb+8FeUOrpo9rrqSWQp/rKd3B/R9MifzsLHZaTMahadc9CRZuMBnCq8C0oJs2wjnU+5emqFgJkV2
mogdpA3MMZOzFxw0NcDsqPoVV0nuzhYNp5Abt4s+pnn0M1/EQE8cUB7pMSXvTtrS3//GGaqkjQ3q
LXsv65jX/2iFIe6LtZEjJgYnY+gAlM3noZ9LzsQQenZ6MaG1opDZCnZy+PZpcYLBOQUSf6M9dQG+
S0JxxAPJE5sR1pwwM+Mx3kC/o6/3QvlFMTXc0ZZvyQbwuKSzw+wHE5T4s4v1yefA/iO0XjCY07CE
QamClM4r+9u2dEUBTyP73wt+p3sqaMbpUYzNJtModitcN+9X93hEunTXoRgfmYduAHt6dMBUi3Ga
`protect end_protected
