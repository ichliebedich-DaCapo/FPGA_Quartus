-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
onp0HGzvC+kvcJthcvtmCaWafJRyrcWXbnUKtpMOH/WQJXTa3fXMCzz5akUusX5hcR6Wdbscay5U
Y+UF5tfTJez6iRTeG9NEqkMS2ruqEf99qPVdqk0v0x+MkcVeI6FxEjYCW9QiI1ZFW5IVeXOaBkaw
C3kjo6xSNi62MxThJD+kxNSffMuqLYJIY0vw8avkPNc/q3/LpUoTe44msZzkYUg100inFDHFmMNQ
RZdl7SWrAFWMX7VQZIin8MRy1zKad6PRQRhkYBHQJor98hE6OGwwtfsGBSg4lQfFp8NQPqPBquVZ
VmR+XZCVk44sP58nzvrCAtkzqx91IwvOx+uecA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9104)
`protect data_block
+jHGr0zsKJKg+xm+IHsw07SSkbh74rNWJtHQWgqNB34l4XJqGk74nNq4xghx8z6+xl7PQoxJKEMp
noeiHhnZ/H5Miy13D6zKaQZ+OIA/P38eOQQYHFKdifMrBsnyD1K+x6WTyrKNPm7vVkrlEoDcGx0J
Rh8oEbA+DOvO4B/i34cpvyR2Fl1T1+VxajtmWdzPIktJy5lD2isVFgXIZQL4ybM3iX46tgT63Gmq
awN5yWdnBHJXjG9cRnm97ovz44/nBswvtyd9yH7o5LUp4Cf0LkXtvXUux9CVWVbYU9qZ3SzsJME1
GTAYm1LU+6CZrq5rZK5eAI99zuUJjazseVEBWC1hBLZIPsU92COj6aw2nab+7EcTHmTzbRCA5xkJ
O4WB0pDjxGDTe31HodHs1LGFOsfDqtYrRWejmxchJHZZzHOB9rR/ms7EvFwvn/F7jgefAgMsfvMq
GTfUW9LRGciTKl9aRCVR3JfAl1aZ0+yEBeyKeISrfqyVtshk+4eRAPr2dMw5I/aGoknm0/nhMxbK
v52x1C3ifAB4TAcyFLx9XWq4m0k1Vc/rfWeBYgsotrPueDn1QUK+qX7imte9qyJgsYXW1KI/n9vW
oq9slwwkarplrZIqshqfzSl6gEHBWNxhvqow4RzgQU/GR17sYiH7j2xSEeAbQh8wVzOmW/dKq9+P
Iv4XxE/h2YnZDwefAezFFobWSwzYBc7lWTOc7j0Ra91sbpxXqQcKXZ2gEMxb/Q1EG5qvS2/YkMWa
BrRspAfDTP0tDV3AxScAGaczFynzi0cTfN60em/YX+zUlKZkRKqEjkBfEQQh063aNmzJzvWQ8Hpe
nUG5k7tZqIjBbNjfQurlH0dq6v2sKTy+iiWU1MTrAsDnd8RYxOqNOw8SP3K5hvwGT89RgYGnYdk5
9pcDa7YtlvxhaFSmlzb1LPy6f3vFDo0oTDcwHrdEwe06QYCeYk2WeWTl8IIoS9nftSL3jyykoGEV
U8TaHxUc6Vmijs8lTDVGShb4HEIsaOJJvFcsPoowxSSZZlEsXnStc4sXV2VdyQMBzeMCHC1qhsGg
iXdpEbU09S1fahsC+6c1vq72xvH60LSOyn67u8ECpWTdFjEhOgpjtYyj54TYXML4RPelMtXbZuTT
s9xfdvumV6r0+ZB0yqgxBRtUmltk4dsahreZZqPyBWgJwdALNGpcnTsGIujb5TKd2U0tmO6e8teF
hGcI7RZ3ZrbNG9KY2Y69Vt1msDzA5pOkfTBpQJuWscUUvvOfis4P932p474fE6VKK1iFz6aIDs2h
VpKinGEkBjKrOUTm5c/nIOL+haR8NOzXVD0AOC7u2apPQiIPEDmkspky1vrp0w7HIGBCwmjzGD4V
YhE+Fh9heIVFp8qpAmahEks0uBv0SXkG7M6c9KjDA4fagb5JiYVb+8MIvzqQLM94uJj14oFtK3fF
+Xj76+07HVG5ZMFGB2av4YrMOUQo5ylySkDEe84i7bsG3BjcKVF0ExJoMhV46bjbs8k3XoPiZfZH
hDHaelEvlezdYynZMwVfa6FpW0GG0RvulQd+JxrbHF2GCcqRde6xkYc7UHadMwxBIvlDCh/iYVYb
Yj+rYk/x3S61txGMu3HTcc+FXpwxXxuRG6itVCtC7SLzwrxuNg+u184fbIbxS5i0sLr6ZQF/q5ty
288qOPIlxgaPOFtTBG3JAGMEYsp2eBWN3nFuYgXXgmMHZfcJFO8IJKxRaj0K9MpuV9pbe7btfehv
SdA3/GtlohtmDcDh5ih3eUXR/l6Doh2dZ3rB13C437vhsKOHCyKLWg4orkttPjYo4CHhzHIXkqFM
q/fY3j4vGAa6M+XtXjOxwiP9+Ke+pfx7ImzVtM//P4KFiVnvtsbUNlFpMq1tX2yOva+uVzqld9DF
krypKMG0A3QxyEa++ulmvoc2ND+mxWSMPGCePEUEofYfTuWnHmRu8awS0DniG8Bs8Vj3hhXvZyaf
tdA2ialoclWqk9WSQ8QO/exNVB5h/lTuLStmV2PUm+7ONXEDv8TfhCTALFcXmgp2Z1yjdHdTe0zc
um/GlZZYKAMpWcU6uD0JoUJG/Z6I64w8/V7Re/GTDp9kaO0uzNKCUyaUeLhX516u01zAimZmj207
8vBBztx+BaYrOjqklPYsA1pVohx0mLujWaoCJu51i8rOS+HXWprJlePkxPiMCbOBmM/h0gK2mCCL
HJw0UmcyefDgEXlyokA3q3viGXP3/arsJ2sTu3JcBPvDFnRR0VuKKjlKtNIyWqJNUr3ADfa2RI4a
BrwIYCIkNIMXdCE0TR81Ee7HyiK5wVCIGmSrd1F6JibXjO7TQPeUlrjHCGa2jwrR+m25ZJhXwjeM
HzR4rrwRxpvDfA5MKlFlSHzjK240XhOCp05W2iPh2Mg5P45sZ3712hs/h3S4+tNMLLHiHKuPvBin
IGQvfswDyOfIfqDNJq2NeIitDm+II+iiVmz0Dl/exsBaCeOOItiwLa2L/TB4gJ3AqiRsL3XxxtHq
QuRn7bKEsg6yLZmShXn21bZyBAS0LIUdUuiZoBVlRty2exsJ9NbvCniKzzMvspCxiNGedK8j9/pd
uZ5iLNfpynxyU8aiTcujg4oJ618UbTVn8r3bfqeGCjjxbzT4ja+EJfVVKikr4nY3C5eVT/hceo16
MlWrsj/unJGp/0ZlIjQtI2fui9p0ubWt4NETl6hhyynv8/sE4F2SuyoH0EzMFhMDswkY5uFKRYWl
M1vPP13J/PTf+1hWvKsGQ/U+Sk3KYWjOqZEK2ViQ0EggUyutqLEp37givrLZr5/NGUcbTu5codXZ
kn8iA9U2jZHoTwc+t511goEn+j8EueJAvlJIMf7FYFASLE7rbwW7+b4d3Ys5YARRJJnfXENFLYsR
ymyfEbphrvhSNeGhRquDOP92wyFal3G0aQnpUliPGp9bDlqh4D/j2n2x36wNm0e0PLm65htIAolC
wrnjdC7RIQm6jSvikT5lxYkLN6dR6ELVZL0nTEEhoT7Ynyndw/BRIcERqzX2pdI0/xTALg75YhLU
4DyAIs2y7oc/yaF1vQAM4M3hwX6XGR6XFhZTannrasydKIwg/ibKVrVD52DP5sycFRFLvZ2HQgvw
JSYQfoBuVRKAJN+GhxNgfS76aJmKs1pZ5NYabcte77kqYhxZb0onDfu9mMiwB/6PBqtjWsFMhl1P
VD1ldapBejsxairsp/nFTWKJhdi5vUDW9XT14JWSJCyEgkzyOF8sTHOeDHw+tMj0Scu/DMLeB28s
EibwEjhJsGWPuukIgk4r3I8INs1hG7+CGdAkyuMHrDLkVYFUb/Hu/T9yE5QJdv8deTzlfOlsHjgu
PasjSqBmNxpfMoqy6us1JQQg0MbAfNFQphuaFzWu6GkKT7noBhFajosfuUgCz5wxE3RztBkynEqI
k3UQtQGQPokbBiEdD5l03qBezZYMI7go0zyzvEBHw5h2lJlpDFGIHr+3FQI5SimRBs+f1/JU+Jf4
3XIFwmpI1hKOl1BhbDPXDiR470twxrISmzcEO4Rdjh4wVKawBGcuHZBPqR8p0gJ0ufRcp+kmZGWo
/EHICP22TGuJgic2Em3N2JwoFZy2QHtyZ8n+5lta7iVC985IhrhbFVTKRP6GEhvsN982kU/EzY1D
YkywHUlEMSf8pFo2vtwblWeAXJgKpkmD+nDLZL+nB0HhhKbC3xU/6t7aW2WkFHAXyL55v/Fb6upR
rq+Q0yvb1r+zY2EIuSGQcrIUSECFEG8SKn7cIWbxdG7kG3DkKGFtugIKrCEFElfsBIoJ2wWhlfST
dzHDNkHATyWU1OjwnNZtZBjNerNDUlPf2zp6UFVv3Tjh0cpxymtPoVfAsBGZ03TD8HWIVbsrE4O3
Pe3EJIyg95X/tzOcXvBPEziwsK7ZT0daLrADi1ho3Z31tf/4KRAIW49cNMN3p8JZdmQCtfkNt8RX
qEPmmHijNvQMwQ6gFuwl4CFM98RJcHrcfNbThxwalQXehsHQEgbkfGTNiIJXja+XIxotJl1ChsJT
Em+E8FsG5bvR6UQP7riKUWiVx8GCwb6m0/HgzXUY9yT8rgZkXuSKiZh7go+lKhle9+k6lWEKyPzW
hPXwFO/GxrevWBZXrQiwUDnj9p04onwT0MUHhQH7cao7bF36g34JETrBoI0UMc7sC2pfyCEcKBGX
nj9zzil8hani/VYG7B0CwT4aOVlcjJamKYRKDQ4L/nhe9tk6PONYFxTYjnewmmJtOoKEZT0CL///
gnh/7IFweGytl/15qyc/8MVf8FSYQyfj6Lr1K9fiixs6ISC91dOCLtTaElRb004ZeQPlm70S0AFj
+1SlORS4Y3McibnXr3MdRpULfkpq37Uihu2IeB71qlfLLws1KtzdqfMtbTb5RYVQjVN5exKeXT2X
t6BdssKuD824ZHP6FDJNkylm4ew8HtQdiqP+zRLmT7KI+HZYzHABV8XKCoXw53p+AuWYgGfv7Zex
XSZaP1F+OK42Ewg7X+pjrObpMmxT6zOfoKJQfHWeHe45EmYO/g7yuJO2JOQQlzfBiHJM3Leso2z8
BW2RjbeQMWIXm3O5yLT8AV5hGITZzYfdMVhMLkC+xStnjKKJUBqVHkINTGvD+AjdpKSCR74wRQx1
nLpJypzZSjMhAdkgmR5gOEnVLOpkOOQpG5aQFBa1uTOiidm9PMgCfjLcNOxrAbmYGGHvKWyfkfSw
+H5Yxqo/3sh3ITNkP40MOGAt+uZRExhpT/yqGfLC8rcjvNE1d5acKG4TLmr3HdpfL3HEzetq4xsv
ZIMG2rmGb2OKT+V1FlX/mEF20MxhK1c4C7+svuIajbIIaZ8ZD4dkIhZWXWB8KdofwjKu+BtES8Ze
gouj4aNmRSBQ6Fvu/I4iaP6I82XuvS5A4HKQ6RYjGmdXxLZphNj/4tOzNqojMVTNlgJjfiLkpdyS
OgoQaH/DxBgj6RKmaFrPF7hiqIwCrfgXkcpRX3572UEQTvvL5be6pUSNocCb2k7AcwS4pICE92U5
ZeI4uzUgMQDw/sdcYosb1SWSR32kjm42ZuIZFJXdUoQ9gkH1ubNuroH7mjqsmY5ywERLdzIk8KbY
OmrLB7+dzQrikVRB0S5rwAOv2WbmqFbnEIEY5LXxdXHyxXk0/vi9CjGVFAp1t73BT2q1WzuKLWbS
Jjrm7M7PxGh5wUsK+XFqudhMKVxvW9ITaVSi/Jg1VbLK8kkel0mlrsInZqyvvZrVNK5pVs3db2S7
JWoFbMxNWm76ZdktRtK32/PVsAw+rrEYuv6VsPBwPRvBMDZcbLIBGZFSIWW7CpxZ06wn0JzFyNce
GnNpEs55bbsofRBMa9I0A+/b7G+44yStd6gdJzgdgPc+vaUO13cQGsxWwD3WhCnDYnUZF52iqWtJ
y6UI3XslYg5ESEDqXNNUa0oRCAsXAnYiEHhnCiZJhEgDSKMG/7aH6ssZw/Bttj3eAovrrCI1eGQ0
A47WZVMms5HWEl9ci5eIBT0r0jExWR552G2q8yk+oGkg4PVpi++HDvP6J/wa8DTh2YyXFNXWpAag
9Oy60UC+Pw74qR4qDsHC6dJtOitEzac5JwQiwnAP5eu0eEDMNGovD/C7oLMPOEzVGs5ibDnLxAkv
LKYxwKMh7jNqteN6TxvPa4qfNMhImGCJFTDSc+amSFlqoRZo43M+ArvxG/BR3gp8c93azsBEklim
X53YhFn3ioTeXsmA2JsNPr5Wm0ZP2/a/ofQKGbFx5+g0l1OH1bKuZnjUGrlyC9/CUpaHOo6TEtbj
fPqGpbW+UsKHgiO7v40n5KSYohlEgeDJTGOaSlPleAokpxqVLjTBd5Sx5Zl2hj7pbUBWvX/16xqQ
A144loagrtnvS9fo4AaH/ygKIMwmCjWVaPqNPDvZBhwUjm951hy2//YIO7eurJcAKr2bYlo2erTY
momdH4/15v0vvenR348L81cAEAAhPFUS/Uy25rndTaAfHyiWArbD+uCGbYVKh7MekPwdkskZbT67
JUKyHPXgR1x0FgxA3H5XUv5egsQbo2gm8xBKNBYSSPuuFxdrIF6+vuibEUDh9t48l3Tm3BEHmtvw
MErXyyJBXgX+ViaO2P1ETzneWNE8m7xCvEZYBMWDUOhItcqHEAJDCe5G2stwVeiUW4YqVo6LGgKr
61yDCVXTlmOfd/QfV8dGbR/hVJa74VpzxNHDk4p26k4Q1PucoXSHE55LGsJYxlmHK5SGCVt+2PDu
l6pjA6z5WVUQRisKWM2UKsqyL1YvSgsNYsULiUonigeYPk20chHs+EHUmSemp5of5VH8gweR/ioZ
TwFgL8PvORnkOJ7HuDODAtm0mQnyFS8hRVShhVtkht4lYsO1AuXqd+L2A/cXHoEGf/LBTa8Mo0WP
u61wKNv44cw4PscXjcLApY0kGqiwQ47eGseRgBU6t4ftADWI/To91ngrf6Vnkrcoq70CDC2eqQ0R
jV5tr0CY4uxHVtkW6pjxCig7bj/IBf5NHh+g/2InJEvyS/I8ZIDVVZKy+njAtIXJJvLxSDuBZkdG
dgXDV2zHZuaLq+4eaNdU0D2XqTR5+wF+DqKUCmbHyxTjWi+nM4GKxoelg/4ATaOBJSKnXG5LkCGB
nnFcQw3Q6xK4udkFe2y92xaugeGWnBN5AVlLHFRTAA11vA4mF5VTtdbvPFY7fZne+rjI+wzG1vd5
48ugXXUcFdTBqYoq7hJZ3he7rWChxxgJyh0JaX2I9uhdYftUCHT5KSLmmHxP4OZYu/FR3IHIt5HW
r2HdGo+jbAUzr636sU712svZmWHB6pJfhjktmWfTCILtxdAhgZlelEXJhYTVFqf74sC+h2RvBZA6
N3tTLFs5TVTht9Qv7nfhQ2ec/Z0yH1hQvkJlOp4D4aojuQFZonRLpQVlj2ibJK5VuISGsovEnZqd
uBNdSTmglY5zHqQBUxvQKHKIE++l1kylPUhDejbgN1uOO3Im5enT3rU/Xi927azrRewz/gUTC1/q
ANIuinOufvDntSCIrZ0UWzG4oZA/crUbcrhCVOk9lsL43jxwGySV6xmitP3uac3DOTTakiBNslf4
7KssbbYiKUYzP2yIek9DA6ycAbn72ZVdwLJRAkX287ewiJgj25ofCbDGjNuTXCB0iKYgIzxxQL+1
o8c5algRIr78/bkg79ztcwDxuhkrGNbMfgnCHNnxXE5VGUuZ6NoQ7heu+vPpK72nURMVMeBRQekd
C/ln337x+WdQV034Sr7JCAxTAXEncwhEmJB5rlXdWuRHgP6eHpkvqAJ5PJl7tunr4k+Oqx4qfPcf
fxfMEDaaYsmVQ1zX+fsvlV49Hiln5gvGnDFzENIlmHHOJCue/wK9L7tijH0U0bcplbFRmLAIFZ0i
ntgIze7RI0g6MXeonwdMeHLdyOQpdX5g5P0NIgLhtyxHn0+jU4Vdceax1gSxhEalcsCJlkKp7ezI
YF9M+c6byNW2wv2b1Vz0U2yQz/8Uw6FNuHJx+GWO37d9Jfw6M/MXcdHqbOud5FgRPXs4vkjX+7/3
zMlA9FpoHANsHnwkokWUcRZDP4p6VvJ1fUn5hOlzwOVWhMELprA4VrXP2bSMMoQGPLta3tTAT4dc
mU5uBfRbLwSitrde7NQRJRCbhY+j2sGNeD9fO8/v+HmOEvmtfupaygKfnqDOme8isPYVtXcHuWPb
5MZJKWj6w3WSp1Ad0bemEDgDuzRirqyMJtNVrh5Awm78xJfRy4eGjPpI5tmh5kU13sWSOvZk5Cqg
6rwdw90QmppbKqQc5igY0vVcBdHbEMpFO7kurGmAnf3V4v6R3W7DvgDs+IvFDLyQ/z+T3dRWEaue
C5ZoJ8QyiepTvZfPq7Hk7BDDY4FQAidIF34tqJYklausvIzC/cSDgxYIwPRs6KqsPQLp39woCXdP
43p4YWOyGJnFNQ929S5Fs3s5roK2DWA694+HaRKdrmjyJiTkGFPAExjXbGSjQooG0pCJS9eIKzg/
mqkgYSWzttW8ZnaCAIlOPMzVp1aoYtdrUpOHlW0XbduBXlGCOkkyGBhwDKbihGABnw9C0vjCkUEP
nDJ5T3RNrlsgXF/thb+fk+vPd4lBvq8uqYmznMNdbZswxGBaIL2o5GV6UYCSTyt1zdR/pj8EJ//k
0unwQle4Y9rPn7WVDWt9LObgLRFc4dS1OlrakAxAlaP3hiMWxD/Y++w32EDwluI7jnqV7UT92LJh
zguVkyMP03DOeM0Xve9yNnJf/YcT7SyIk3ZtbwUu2bRqVlX98gkU+XqJTgQbXXAiNR1t8QqQlI+Y
pcbmUJj6Xs5KG/5BlJdXkR99xPekY0fi8oaX8DoRygvKojM8Ftj7mdHEWzj0/qvvj5NMXlWALEUM
WPWG+TKZZrbk/KiOFhITNRPc2n3mCdxAnF2meiZGBxNpsA5GkwrxifZq/LLXpP61NGFtXTUSVL8U
YskhIpIihIFI5jZqq1I8QGKgLW+umaXSa582uZb5S80AzXhFFS+RDlDIZ6FAbdTOeT4fq9Yd9e/g
OSZt9aHjq5pZ/yEhYTdebrVD+Iu1xMXNs+iz5AB/Qmtc+Nc3rWi4kdyHW0xgCa3BjJpsPhQJ78/b
rlg2mywcRPBE8wyDjVPw6FCMQd6y5Q0EbKQjos/EHquT1iXR720ahxCFIenfNBpTgavfF1HJSWjL
2vZcXf7otEHeiyD0cP64ph1UwBb7A1ffSn5OL4mux0Jgg1eZPUNJnJFEEs1lehzUarnmBYzJL+iG
pc02KgQCecFMyIqHJofzkiNf0N5wn0EH5kA6j59rtw1oczWdQNXsMKoyszphqm7En+BHeZCAsTrn
loroizUWvOJTT1bIr4FDk0ovaYVaXh6R1auuS4O6jThE14zRj4+VECaz2sBVzvDQVJE8qYqlLnUq
2vd3VQWGyIjEmtJ+Jmd9KqLElj/cY5J1uuluEj+i6Omlfboas08klIyrfZAwZwq6NsEP4KrzOghV
EW3MZJpIz/JFmh76W6sSEJkWEVsDQDbMUOlhIkWRCzOffaW1CrXtaC5zRFFofN8Glr2bk5iPmVP3
gxR1QPX4zpc61PJNb7Y4vpDQ5O1KjrLqQDZiBWJ/l56fp91YGAUdMatAkEAu1QuNS5iE2gYMjas7
+UUzGWZn1RfC7JDSxSX3PbD06bTJP8k9YOl082k7ViACnBbnpZWhlga3xRfNdSekQcVOZ3JLpMFM
Yqk6iDKJVT7E6INEBaN4SzaJWFTklvjjFrBJ9SSuRhbR8EKCqdcygqOEwzW5ED2TW4Y9vY1lX6Cj
cThP5gLXGwZRPi4ISxr+EgjAPjqSAhuVueOysUrbgHt3oaBUuHNYN1hFfw5DdppDO87uHBxG6hqr
Lg9WRsaBe0sN6O2Kl9PFVn0EmsP8xXKpEBB8evWOqhikExB18BuZmC7W66PojdVuD2jGud+RxUel
BjG9jUJabNdLJPMCzKrZjPSe2DAu+jsWLQhyYjpr+foa1uK0whdkbYDQ/PnxXITJwStJCt4G8b44
g+QDa0hrudqwkHM4HfaAcUGxm5/YAXYV2y3/mxQ5pxaBJgXNXYb6OiBJzGgX1c5rl+aDiVEPs5IV
uAlH9xzHRzNjFKfhfcxURdg9XoXfSaNk91USvG1b/wU3yW4Fcjsu+7PZhx5jrvub+zjDy/98QSRA
0oAJ7Obw+pQe97rYbdILKppBfemMayIpSxS3lKDQ0p/Ck1VZ5pS7ADbIxSLOYIZqhUYDn5gWmhaT
xs8nwZbM7iJwkqY+dIYRKY3i1itVGXraoqPVbA1Q1P7VJC8aeZIiBGdxI35XAF75ltXaFK56Y11d
uWoyJ+EfG/fi9qctbru1i/ie0wGG0odpG2kU7qygTs9ImgB0fPK6hNL4rZYg2+aIcWMmayMLjNfh
1SPkGN1rg7q711DFR0sOU1XZNGKTPZJUy/1auZ4OgWm92CsrwSKoPTrUibf03mDO07S5kVbIHFcO
7ddyVrnIuYzbEm5x5V/vOKpcQiWGvomwmJ3XbLdUPQntiidoJ4WBSys40kZfbiDMPHW6iSHz1L7O
nUL/Itsf8zXvzJcOWEbdU7bb2KmVOsSSLCSZ79exythIsYN9aMOlaKiPEaYVJ4/ZxY4I+/Z4JEeJ
M15/IrUfodqnhfMmgMqUHtNobvXN+I9heU08r03l+gnyp8Cevm3Kdgf3bkPLOdcAtb9U2NhIiHUk
PgO3kXkWc8vBCmTAY4A79fnu9CSGItbg5i5XEUg8/QcTpdHZ3BHmmtS+3KLRjId+H+McPz/sJg/t
SiOIUEVbUjGi5vy92M/2KIzNTtELwsOXlJmMT5his218MOQYbUFZ1BRsp3yphYCG6rcR7GFV9RB9
nd3oVVGvruSXLKtppC5oU+WAciO2YERhoTLws6OkhNCwWmRoAqBMcHcxt/OnBMgNe7F0eAE53p31
6FPUZJ04u1ENGxksNRtDQELRzsjZaM++gJJuGyp8IkyPCoQPqUZCpGRz7csDoA+1DoZfQMFT0jFN
07AIB7pMO4wwy9ExOqhnJNnKun3dyHvyelgmlu511Rs0elIXO051e/6QPDb0L02p1fk8zb5DdI1o
hWikfF1E3+8xStgzyEt0qB0IVuVnN05HXNzlO2Oc9Jg4LZQ2GfFHwZCp7lz0DJAxzeRFockDTl1z
p3WcZISj4Q/bR6Bd+tN0M/2Kb52yO8DazwNhg45+V6RUZ/Y65xqeENHDS32EwKoFskxHlE5rdCyC
VTUcCLB0UcINb+Z2BkZtCUxr/G9UdnfgMk8gOgc/nAt70Y8+fC2woEEp2UAuAfXXQYIGwQry0rTm
KU+KOYQCYCJ1UegArir1WscmZqSd0sIXREkWfgwpr0fLxflLKqmJIrxy1kZQsDOjAj1jxrPuSGoI
2xymHNzMy4xI/SZZ9xrl5/M7BEUGPHOaTodIzb79lpz1A14VLKsbUm0pKLSqWOTFLld2ERAoaDJM
+PhGto7FbYQY158KVnyDFIcvmdsa2h6lwoNtBiY5/yre1LxbOv3QwDS0JeZPHLFg/gzjL8tOAmnN
C9s8leWyn3NXnDfHDdB1W1Kq1wlAuzyDFaSEtBdRxVtIp4npAnsYTMBMEzkH46VnDU/oi35GppdW
b93OqpSwGZ4IwfPtesfhlu1nkHmQF7ffUd33nnHvvxFsZFyntZKZBv1C6eu7qpcSieuDvfyNzmmA
M6tq5h53M8gMEXlMhC0uwiFoo4IxaFW+VTV3GtzGjvThp5Vn4n/axkeGGKPbO8mt0M1YFMlIM+IT
rZcqeyOjMRP9A6t+5kok/ONETRpzMo8YBI+55pTXFiE2e2ir5TB7RCgto1eRZ1P30pTbn+1G3iJQ
w+ZMp+NEPmQT/eoolC7uPNV9xbLl7xl6LJC7moFbjdnmq1cKIPDh6n0Ki0d1dIqx7uB10iCgiMUP
CW7TywnpNX9y+xhQg8j6L+6A1UDNMF/sRUMozZQYJFy5Qy/6VEulQnOkfjqhKvGblvrNf5Wbv+k0
NmdQxO1l8AOji2bMsRYlcBxX3GMUTfKbvPq+8X0rSuK7czihX7kO8RAjVJe3HMJ+uA331UF4BX6J
dMXLLnCoW1/8/0ILSpIvlTpOoxyaOrtUBJD9DkQjq7csJxfzkunThu9S+usMOJ4JC//kg4/rNlNY
PrH65brx+NIlyRi6V9JA5rypxS5yd08veVjnh5qaSZDx9EeTjubiuuzP1GJmGOYo0MRKrlNUfv6A
1KfQWs0qeQjNy2rbeW79S4Wl1/SfUAACKSMaR6KyZBC7ELsA2vf5EzSC3bESl5E7mhFd380TYhoT
qfYGjHOjYVqoibb7Pvp9tapTMFLDvxXdHUfK3b9TrkwxV9bwoLxI80aLp30P/Zgk0cEP6g4HnxuM
Q7dqfbx3pm8WIEBwvPmy6fRsXDTVqtnKi5hUKdopZk/zQQMy3ca+Ujdd93cnkXa9P+HsP2TgNarz
JKGdaS1oO73quAdYvaP5Hi2AHq3Xv2Uw5KYcYLde7XzHeNas09efRLvOkfER9xv8UKOgPiIwpevY
DfB+5NV6y/hZCW8UKGSoojJ8vuDoAHVr19gC+2pe2FelT2LNLkdFqOjRQpPcH5QA9a+BrdLTxBCY
ieQcOj0RTOJWKX0QtYjwtME4fUl7UoJq4l42ZTsZsflPEHFb27upLLk=
`protect end_protected
