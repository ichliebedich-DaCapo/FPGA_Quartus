-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Z03Nv/mTxKA5pPJITTVN0C2aCMuDF5sNewEJ5EDiHIA8t3DHHOPXD1DTKsY860wRSneRUNJYB5TO
AwXMjbQzQaYBGmB9d88WOSmk45qilfcOpSAywSnLk5a61v1uHWEefpY0voMAiwjDMLIGPBF2LZuq
gXbcnX5mmpyNZ6SiuynHVdfAWyMjNV+RD23h6LvU2aApps5C/gIy9oV3kQkYbxCF7HVf8pnzRHjp
D73VJg1IR7pl+Rvf08EFjWb/7ORPxlIhlCjYcs6msJOdFym+Aes/R2B8X/elfnWyaRLIzoOriHm3
bWyfSWNzjmQVy0+jOeL4FVCkgZRE3nKEfdl4Cg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13616)
`protect data_block
kDz2V6JcZ/VoLvMN1e+ph4bX9AhPvJ0bnzmM1j35bwu9bg1Qo9/8i4HT5O/LnArtNU1VOYtrrBYF
OjLpJ9SmD16Kl28VF+wO9/uBs94Wmoh8pu0gux5ZnLCBhN/9y+1bI0PC7zX1D8VifwrFWPE2erF9
1rvg6xQ/z8qhvkxb+qcX54gcsmUgOJqbmKvsxSrBxABj0mX7y4qbu3TYbTsyZLRZyAPgvBo+wOoy
ELHHiReVNPE3DqJBZc1EDnBWgg+mNbnOK40lV/bOHUsJrcNE1dPorTQeKdh5Ct9dTE9V4eQq4JMy
+z9DDNmkMeAeu4SoJB8YbSTRzHoS1oHq3mmhbws2NHdSMnGuDwxi4niyLw9ZMeZ7rTwXNRIEClA5
0jsQrkpX3n0sZMQdtdQuTgJHzG8g4xe+XNcskSzOFiDRIf7zy8QHHCMo4hqpJU/T/oBVUi5bUw1W
B2irr/+lcC0Iiy11axjij9dRfrwUjYijI89U20XHg9Arv3VfwIYvbxKghPKvMtoJ4gcKnaiBd2Y3
yIWTyucp9N08X/eLGcDj36JGagBKomgn21wgbQmwr8gbbMMOhvjApPQ0MBt10nXt4StH2GnntcO3
KratGgK8tJYJOcZml7OfdzB77IFO1dgHHEvI0lXhcFtOvJ+qYjJ9GN7nC0aPNs9Rtw6X34tQjq7k
WuAH3klPK7sj8XwsbUrZG9Mg47Pyx7rKOb3xn2gYOHZqQ/3rf9Sy+Xl8adbissgT/vT72ZHk2rFk
6Xx1W/IDqfAVJkA01esu7+HN9vhUsxgqx8qM9wxzfIaX4we/PgMWQgCus1+6IQpkIwGTOyv6J8oy
1L6RRSFqhJw0dWgWExTEoOtDs36nGJvvuUCWXDqjaTZ3rOsaS5eJOBJRds7KRBbrLh2/3R7xqLNH
IkDp+P/LtopdNjpTQY3nMPGBwckpOIiw1FzZpfpWTu/NPsXFoKI88ltvFUoVeGPnjGtNFXWz0xB5
8I116H1e9w6NG0Vcxe3bZUMSxXpCKrgl4FMyb5ZNyFLjEIzuMzp8F5/os1drZNDh6vnvffW8xcmX
KDrLVZ2XPagbvTkB1dIB0qLMoZu2yIxTBxYcXzpXETEDuZBIqOIgj8mh6UFsGM3mTyByHaDRKI1S
9dLhUlyMP4k3BpXmZ2LS7kkkh3LBZFJL8TnXzr3X9x6T6cuT/GAkQSneg8blIyMKafaJOyRVRG+l
IWDyz77oApriIQ4yj3tZHiaIdOl6pqfYNGQ4DBc2MUNAW6l1SQeRb4yueO0Rn+nHulyryg0ScPOD
H4mDgwv5uvv9GGjln9co9Da08yudYQi56E+TxrgHDwB9tfbAFPOSG/WWgyL0YHbtgoYn9pIpOKYy
BKxAYpw4y3mGrPz6QupJ7fSk1EbXaUl8kgEy7lMzmFcjlCVWjmpLDs/Tcjbjq4j8HqrYnAQsTjSt
uWQJSeVi11bQtIau/vcNvpHQFahKdZYGhax5bGMkyVj9TvKFsYrcApSMoRVKSWAwdWFRswkNVO0c
SrdyBr13ssnYR08eY4d3f+/Ld1R+tD+eWOmoLbPGvaa9UaBvG3JLYmNXw9Y3K9LKrkABW7krXbAw
EomNG27yf+5q0ny8s5rjzcHcPdi8yhtdiulL6Qc27LF9xMSQT0AVmylNj3xTCGtzWUi+Yi9s5Eay
MIynRN1slrk5XSPesv6twciOLuncoKEwRDgb84EoOtJzCmGyFiVtFjCdbmLERhJ1S4tlykJlwp8a
h7TjzlNRkcoCxoCRAdwlfsgnEQdoRLT2PYXS2+u0ihgH3NFK4pQY5tgg2g5QDUJi8uDuj95xr2Mn
BAqGoel27Zh+hVbsNtz9XDYiZmuTTXof62qm825vJ6Hpsa2g+v0LtksECzr+yDofzwArleh+8S/X
c7CRsQl5tP+O/IwvTWBNaJ7aq2aa56yiXaemadDF0AIsKXppJ8WFZqF0sPgcIAfWa34WAbd2vQuf
B62frgh0bjYBkHPi3PjkC8XwFm3baf+TmbHrsT0SMX2JWvtd3jFNxAugDVqZpg0WxG7leWPkMsFl
zQTxLlMcya22JnTJaUq3rAaF+HBh67OmjoWgsIZ7WF3NAcvWK1gS1XEgmL7TsXfbz87d4WILHu/S
U5fq/1b+LfgbvNKXzP2jIY3VyATJOws/d2gZ5uVkw+dYq6dYnIG8RaY94Neu2rwnmYWWKT6pZgxo
gHZY9Q9nAQxPUdcgOwQOWAZQM9tEzs2+/MsAYQJ0M4B7EbX7Cin+BL1+TrMl/hnGzVORqvjaPG2E
0EXrC2yibXtMSSLSafv1ak5exfUEAmYwp9T9t5P75TcR5dqHDuIyZPw+W3xOAD5NhL2fN7RNuLFQ
5ViHqVGf8+gzDDds4r127UXnkriTgLB056lY30UIgE40qTVq7d4Dq1GxEu49+ubqEXsfxvIVh/U4
iGEadsARsM+tjVAsR2NZnUBBN9hirkAMn3KraygH1sUOhNeF8yY3Wquvy4BVMJPnDLi/uUGalI9b
P+djTe47dy7KzxAoF6BXtV2jeTMc+4Oy7Bparkjsy6L1E1PS+AjSirOOyEqi2b9GoInGC2SdaDWY
W64LavyAJtz+OhMH6NostlPZvYptQLqOcDCScnpxnjGg/TLk/ujt9s5WLTzYNMk5D3EQYHK4/O9f
wYbi9v8K5K3eSTThLcuyvgVVd9PJxKV8PL0xHEr+fachw3JTrV0D0Kgiu1E70FcdQepCebK8mxMg
Hi1hKky/fmBL3YZzgx3Up+YDux43KuGLEn9Kfl1IbgXZfKaTQwfMfLF91HwnInJSIbWTaN6DR8S9
7CSlbk5gwIOywqhvRn0N+AWJoz5ZTCiqrX/mQcjtftxV6vwRDQ84UnuBqHwvX0SFqIhGS+4eR0HI
M7tfjxVdBM/lv/ZQ1gIkdj34xTJ6mRsIh+qcEzjeqsgHDe2zWBdgeTY5VP7WLd0bOVNrmnVOqNAn
Zae6M58U/WVZ3K4J1sU4sbDcZAv7c9d00YRJEWtaHtvd8T6TutyMQJxlmtmUeBAf9WYgGpNQEVUK
F3BId7vPcxIpyxzcrvFbRFYMX7PmQVgXIuKXc1uK/8oZPCdkKT+2UX+Ep74xEOpONDR66tpb1uqz
m7P30599dqc3RENKExN/taD+05VcFcX3vL/Tzc13pjR9j01WBfpUimG0RJofrQWWU8wBvQYlfNra
5P+eFPUnLg7UuD5aLmamqf72REcKkFhpiZxXyn54qWZFcfscscQM+7SUnmh9l/amxzikq8fOB9XT
A8frGGuR+T06Po86OUX4d8J6ICgQm51i7YCGhAusQpcmvioORC3yRDQzXD3D6XRCjymeR0gMdqA+
4oWjcTzxNDlaxhrqVI82/jE3vEtpzlToC4hs6jRVdp3LYXkeqQzdIzyF4p+81ymfboBzRm3U7Q4u
oVPcMXwWJfaNEqQC14r/jMVsHZOTzVwZEh32hHFlkvG/deey1jESmPUw5oBGoxXDXe/XTviNJRxb
Iiq1AU8ZXhHt0eE/mPytE3ztz5/6wS+ojFMyEsPyvOuXNO+17+TymNBVy8YZeLSEibBuI64lBBhO
cdFssAb1dcNNY3VBDDV0xLEpWH/GI20+1BJe46090h6EeWDWNoC/pwdMf/BCQEcTrnlCa2S1/xxh
B//izJiKfzYyU7cmZsGdp6r03AipEK1vBJJ+0GWtbrSvsQ0YyhW1LCIuyy/jxKA0VQVI04oVlfs7
2vXJca60sh9e1LsGDAsfLbQUPEiScsjN5qukyFXd1WEt1IZs5AcKynXd83yhoAh+tOaOgIiCZTcY
ROVWCTot3JPylPTsz6U82dP4FN4MPd1WLKqvWQuCiZfrT8P13obUrUM83hBvJPnnwgybxOBhJCd6
En35nP1KX5zwkp26LTeM9CBCsV0/u37oErv+5lFrNR1ETmslSdbOryHhXXlUw8HTwxk3k8SgU2XO
OGXiGaBglZBW/qzqYkkXsv+cJX0gJcxwsQa2OW9nZCkDCzfnF0/1Citu9miQdCiWY7zVVw3AVkMa
ZUWcizEQzTKSeKSdHa9zC04CHyFMDCuWugB/1DctwldGlGTCLlTgTRdNE2EcPXk29gfndZOsAv1O
DMqpyjwrA9xXifXcNysTd3ZxIzLPIIrfVNMO9yVIm4m/ofdURwm/LDEAMlCZ9g57XrXhwcFizzrd
u9VQdMKRsczDvwv+DaD/MKv8u0wNNjjr6T4IRaD8QV5QXppzk+FD01CZ8cY2amVbPwnNx4NlPOwv
heinZJk2IcKfGGFZhI7TQx6+dVbll4D2uZ1ssidVQINjzhlCsh5qRFuZiMKCI4tNtUkFytDXSqzh
x2Rg3ys0V3fB9ZYzbMT8e6+3FXJVPtMHuvrtthqg3fpyXl1S/RmnR8S0EGEFguwH7I1rboujUUcG
jrWqLVcG06PF0f2TO15lGbyyF6K3meCbxlimVYaYvlPBtFHBiaoFb0uSQKgcR6gtDf1TFmQ0vLla
wvkEiDKOok+HNXimpdc09O/CYXs+0fjaN6smfO+ax7EWbLBzOVH1MrU6YQog3aY4moiBO8prXCV7
HiTqrACq/X7WjoF2vyAFHpoAA994Yuxzr2mV53hvwmJM4OHHS6zxKhaRrs0KaeLRew25IpZDIj9y
FHfFzoAJM+Zgv1Dp/lpUUnLpw6643h9UWssjE6LgigCh2I9snX0fKLHW1BlU7tHa/F/m3XZR87Gf
pRpJdfHwdwerHiElN2cKIw9wXCrCramqj8LAlQtqS1Fb1BqM+MYA+Lh5J1pLl+bvid1obj0Qlsnu
p0RYDVLcUsPPqR4RvEMGUQ6ZHKMRKJvrYbqAk8zAgbiM+AakdrYmL1bnZnjHdlqeUkoMY5K9kLLs
8voGJC43hzM0xL2r6+ryVy2KCdL0V+8oYHDTM8s7ekhPEtQLadS84mmZnZ4RghiIvJIEQzhOeHkQ
tx9c7y7bQv7xLA9wWKH/RzPhqFfQ1CuW55YSokwM6kE58pPx8tJ8r1ehssYmS0L78nx1+5tl2uvf
WHifeFrzyHk+llF+tVTDK45Sx6a3SDBegNqsEM/7xgMw2wnBbiUNhdPThIuTtw7gSy70vG++GsX4
mxO4MhYNz0eZ9XeJwGwJchNhXFIcXhvZ8S9z+BLgTVYUHZgzIjoku51OBXZhcDVYbaRoaNxbmE1l
j6tuCIBET1Utuz+gizsYRz2EOX78birbDCWCnGDAsgqvG66OytkeUptA6nTeNQGNuiTAtUHnHTeX
ogo5s2v3vNznIdcVuVnPjlhHkydaFTitYtCK+ZyAhYD90cWv/Wsx83Nb2sUv1AaLklhURQu6tSR1
3PGA1OZLuGXgFTHBavrjiAKfblbsjuLp0A32143xyyF6rh4Yrw0EyDXMvO7i2ckvFqgHChNUwDdy
vVTSn4tOX/tH2aUo/6/4/OrI66kHuz7dLkKvpepU5IrqU5ERdotT27L03onKGQjOyY/LbLPADvXg
6/n2IpVwyFdImRZbj/0PYeuazJfgg3/6USlQeSp6QfKmNA++pVrUSdLoZGNcxqWpKfvL97r2B0A/
QfSP5Wz4JKaSurbW8K7k14HmZEFn5ezQjpIWFzDYMEc7rcPuqQxsy4GvoasJWzOkZFj1/WCjaOyV
tvrXbIx885R3sRGlS3KFRgRg+kSzzsnzOWjibME9Wg31hN9PyoC5qlBIzmoB2mJnMIQ1lKAWXP5Q
tooNZcEZQGOFch9KbaaJGJvOTFvgjJ50WHyKa6gDujkXNRZtMoYfB2usvn/8cxWdhiIAg3MH0Pzy
baT1DDortqABXHukSwfcLSNhX/IySYVD4qmCaPvrW2DAFFxUe3PTg6Q3nTnY5xOxxxRUQG9Ifa9O
wOWri4K6MbPYQwnSoKx1rXEEdA5PhEFfcN7qGOPxUExiqEXqLElrKiuD4HfKlzPV2yP94AHqRzHC
Nob+rXr+welNO+peIzaZMZyDvb7mcOeyd90Pw+Et4jrIwkqQ3mmNkezFqmlfauCpmRJubel/p7uc
aMXO84GxUs8ZBXqKyZxYjc7vvo8wkmEiO1N8j5UfjyzY0pwHE8CbE6Eesh9CaO4O0WhGrluP9Um+
sqBHGyOTsMuzBf42mjAqUrX0fjB7aiVjNs8Wrnyn7GJqRTUPHCI8bglMrbC2sbsnyuL7WGMbQG9n
FmvaZSpUGYAWFO+58mOKG1xxyUQImptIM7bTDzbtZONmKOpVESZNAjOL8ooy5YdggjgDgxL8g8OB
LupMb/S1oxh+Obotq9IyZiMt3oSHuoC9oWLbTj+va8UfQf2xCcOMILIOf0QlePxsJ4kdNoCGk+61
+aVHG5vf4ddXJnAleU83dfz2y2+9cSyg7jkQUaJV2xEpwH0i38M6wYWk8eghzPFb8K9sgb7V7HGr
FRfJqx53oMsecMOZ+Z5VfGlGxkLQM9106rJ8nlymhNOVyrAVre+Be9rqO4UlOOp0eWUsa5TcX9Xv
QCtd0wfLg2E+kDbWvAOkFZiZehxwlf6lFLTljjtgS7g2svpJQ0Z6F4xCQWzc8B3+H7GnqrvMX2ve
XJdRaZKvsdKk4LQuIDkWmU/Y6Njj3in8/LyUUWcbpfPVCTCWtzzRZsSUV2+g1aCDyxdVgoyrhmNe
i8MZCUFj0yMOe8yntLe31Tm76FO0NBegZ78ygwDWXZ8+QfXHwF8YqjQ0UBTCpi9z1d0gvjrNFOK/
yh6GGCnUCjRzyHKOZZ/MrLGOt9fAOZx49bNw7JagpJwus4p3o+GzLabETcasvL07MQOYmAuUo/RE
F1rz1zuwwg3zHxsO2Df4MgKn6rFFippvcGeTPBgaAMCEcFF699p4hggRQYG/02ACcenCTL/B9Jbu
rOkK9Rf8FyDmMmEV5PIDfby3oIP+DFNvhPC90T3zzUnt1XrXgENL//UHCN1rmm8W2Cf5bZo78hU/
xmpKbUxcQju/A7LCq7j3WIXefG/XIogq3Vc0uODC0flyF9oZTVf+sbxiF9XmbTlPqF/U7Q6Obql4
fOTnnHOMglDRjpMo3BkTjlWvgJSqDZn+OXvnRTw7CRsZ355T4O8Ha1oy6AflPV7JwDKDuSKCqZ7Q
olVL60ljNAv5PqrqE4PZR2s8H3A2pajK2nfviH1ypQT523kOxeRev+TI4XPWMLSeO5HCj0DxMyXs
s+HgG7cW9Sxw5g9VF6xB7yROnETrGTrslFIdpM2MjgBv9KgPb0PCwOA0rgiBwIX/7t4QQVCFQ1Dm
ez4fTdXoqD25BcUyib3FWUtiNIjkgVvDzvZh4f3EiaPl8osaIkZdB/1ZbOuzJMeLRUk3ZMZ/yrK/
3/eZURGDWovGvcbHr0N1kMUi1eRAtOvZag5vBA8ped6OPWAYUEmXrFEI+jjcSMD9RRTEZ1aOZrWz
I6cLjFXIjxlgDsjGjM+e4fwfyaMRtmyWnsWXJi+xnIMUcuznxDwo540NFFkcSYuHishlvoPCOcQR
fna+JKNViXChZtRITpfcvcAGE3evqOuO6afHvA3nrzyBaxokPGfhQJeWBo5J8tGgyDSl1X0Vez9O
vtbJt2PgvoUPJmQ43UxXwYwUZB9+ICltoomrMebD8OzywhAxfkOJulLfWOlsTLQMbppgvMjy/iGM
vmsurt1DLBU4YyuaPxD38UxbgU8zci2Q/JXA0vkPjsK3+K8snyX1t74CgUN2ByZsWO2pVWu4+tJL
IHjVkroqYKVBIi9AKlTLKfXZxuV7dfWurpVb0882Y4n7RRTGi+xeLpGBTmE6FYjx0iTojs6tM8fB
1p0RrcJkb7zwTChVawyw7Z+jH2qyViHD10MchNPJBlxiAYVL9ttyFU8T4s/7cK9zFIGn4F0WJ79g
3eocLhMdMuMZ02T5w06edC8fJXT6vWoASh3L+jKote8cntL1xF2KHOr5IIOpVvgmtIb95FYXnzSr
uVVAPzeKNLYpZVJylCR14PYVdxAq96VnTRL12rNH2ALu9Scwcz8H8shIL3a6diC/Sdumnyg4crYF
5Sy02wEsrXTBa//QBO2+TFfzR3FQXALcikpj0IU3hXMw9+qUZjpGct6CCPz+0rTuDQCFcCGWEEA6
dHSkabAC+sVGAhd5TvnyknxH3HTmsEkXbxTYTZf6daMVGt649qo7sgYHIGoIXEqPdtx0Y7pSHId0
o+mBYfQ5gaekCIJ0+l3AwL5W1rI6myaOhw40TSYwebdkkwTifShy4Py9TMmFzn9cTyGYhyVGdbvx
miR0CEftIoXL0XhhT5z9oT1kiOtYQLxEOx2EshVrNHor2VqqLrXztdKEKYN5VmqjY4kkEms9z/12
iXNi6e1JF8RH8tr8skclfQTK2/NuOkDOkkSTrN0jcKuTz2VyGh693C/OzmcAk4IYPu5O6wZSnYr1
ZZIqgr/bOkXUhMz/gs8d9Do9l8FTl68ty8zcAd9/0rq3O5tUt+yvElZ8DBQa+wbcj/tz1i+4IlSy
kdMN0VWcNEPTAv0xQI+Tk/YgITBvs9ZTbv7GiuHQ+Xzp9jyMIqO+gqtQCplgR+zkbsJSe4KZrKGy
GD7yMz4X7ipMksoNpD9rgpr5U4IM9nmtdKFPf4S15rQoDLHzfTh+DJGhaPbWqkd0dJn9a9I/a6WD
iSa23Gp2hhGs2xl0yLhsEJrS91bVuEDKYDL4PNa6zmlydjjCz4mpIBlazm2Lkp4zhKIvZ3WafUOb
wk+1/v6o18DphAAf4eM81mgINge7bm7fxxDX4X/LPxRYYaYWuGQ8LAo24fQ7UcWf2+mYOPsv7RcP
r2ctUnKc05obMFDEObUIAOV1ws2Pq0ZA6vv258P44jIZlH3n6I/kMJOmbNlrcHlxb5m7kfQi3Pap
2018TRRpfuTOlMJd/FB6+W6k2l5YmhrtU0qbOcb27o220Z6ozbSuCv/4LAOzYfEbdXXftPs20AKk
DNps2dfelW3acqtVrv+sI28m7QFgFBLhpsBqXSJ585waX8ZpeyKNich+g1DiNIPqkVafXpvUXBIL
qj4pflWw8eAHcmImJAkbFoNlo5JEM/K44MukS0vQsTvkGDE54jOO3TJx6trJVLE1E3+9XaEgtojL
alP3zMQllUBFBG+VFNjw4mumX0ryBYtnk4mbUQ4rS43AQHmLJCE+1jyQbvhEYtDirXYRcisybYNk
e3jVhQkdb5+bUyy7hWCmm2QVqz5Lh3ZLMn2w8L6k67d4xFKBTuosofvqKRFUB8vrEfuJzjEeBIzf
De/Tu3SbQT92pLLEnKa+E3lRENXL1HcQEleROJ1NYqw8LE3a86rh/ikOEYYeaN/urCQmGIOzbppK
aU4FOle9ypwbiMp/Zs7VpLeztTNPQjCvCf5iHLyocKklVtJNonPcg880fyTZu2mT08xvbeHnYedu
yVJwKlpoFRfqVr5sV4t/9Fdxm7CZtgMxv7YoB7dTtYGui05+anoX6/JmpZ/oj2d/6L0lziA24wEF
GbEEACjHja+sXuFEIuMul5IUGHFxfemzvi0jLRkPyV7Hv/GvCyNcT7YyzkejiPgyiWQeaw2uPAXT
s3I7kiWpuuMRu7n9bHsfL5uhF/I6rjKO9/Vr6go8r/o9RJZ+ZHUVh2P18q+XMOiu4Gx774QZ416U
uCLt59GjodDNHKu1EYWv+xMb0AIlM7hDfkzP9OiS2X2xgTjvF6rIDiOcg4V5jzYTYLgo9WupBL9q
PQ5PjJVpuJxhXIGEb58nVBb2fc2PL+F1ShAYB22wPTaPGp6HpRHjUWLrgmxfcnlE2M4S4E8tK4Rb
/aVBWyRXgMbh1dvM7CP38YhEfZapcROKdH3YaEVaS5F9WnvvQ8TUQ5j3KKxIZCy9g7dVPVAZtlds
1/F0Mz1ul9Tp8EVwqGGtACl+m3EXlny+dK/Wabpkd0Eh7B/M9RfSZVRThoUm+Vg2S1OyZI+So6NW
qfRU1JyqPpjIYWNqMH49KTc5ebuZAScQtXcykq+9Av8JHhvwlbL3Jwh50uQ2uPwcgIq8vtg2i+YR
jMPTKy68rfNAr3+GcULEV+ugiWf6aA/0nM7WwJ9NxAR86TM68Gpxy6nxxBGXJRxWDQbdMCez04ro
CgNaUh6gcNQ0zBfJXNNhoqLHzpZhfe1rTJuCEWvDdn8TFeG+I43fmwmPx7TT9xRe7QwrHBHdrJqP
x7YUF3eVZt3KAs+cE7TNxqaSf8d7dNSbal9rRgoBpk8Qgzc20hh/7+NuL8AefFAZUPCNyUYUGNzT
diSy4GWpmlrOW4XFpJjHlLdKwCnPxZevwAotuNKx+AmnJTfQY0edy0pcesYcpsTyLab0T4xodSlM
g2GGrVRMqTzNg7W6d8gf4wl95vivZi6GFFwm+yukQ3+CYOR7KPX17dPpbxby5QMlUXjOIygeGX7H
N8vsqVeOZxlZo8dGKwVI3ZVs4o5I8NEdeHJEhb9b82LAhTtYgRbYG93Jfpud5oPLVBCH8l4JckRY
nFQNN1Ft3t8ntBc/D3nx8mUqc83TqQELSYCdXhXV9JTokFBijHZwPojxilYINlQNZEzbzp7p5ihs
H2tY4uUplDO1mpixRyIgtPeHi0aK93BjZ6TFSjo3gmN77vK/YdRBVbabzFbNwRkLn62dy4UojcUE
arYJ46V6IMzJOB3YUwPR+ETxba1Q+4s+LxRmbu1hUHPCdsdpI5QNVvHX1KhB2KdMDRwFOOKiclCd
C9X9zINokWJXJgL5H7U5hZr9Lhw6kuaW1j3fvQQF8YLymKrDnzg2hgckOSCr11yrQFUeb9Vwie0F
kvIMcY036hJV5Wzo48C+jAHZyX4+ADfFoctU3Aakg/SBsowBlb1CckBOh1PCe3+ThuKwxzBzEoF1
M9dh/490QzOdyaex3F78gzAv3ZTW/cnL4mJyox3xQvrrd1/SAtRFpY+ZkFA4ET6FeXuBRjXaQ8Sz
O0/ixqcULxfDyAwf6rUHc9FvVarE+klB7pNyU/YyqcIILV2l+/TKSeVPKCe4yLd8UJ+7i/YujMIS
ASlyJQTOsZ2dtsggREA/mADaOSajk1StYf9LpaARccVUmrHY599mUriZCXuVb6riMm4zKD0E2xOL
Di2a7EJq3m/tIaCJY6W4wwbuTztXRMcWx9a2SP/q8sEiag32XKs/J8hvni9oR/+4+LVC57vlLvUK
9HitclxIL8KTZsjYqb8tp9u+oWA/2bcxaxXr9mdeZdm/RhSPsUaoaucOd77k3Vbw45dECY0Fgkuv
UAvPpUq5/axWUUWhTnBqieaE14hDXe+Ss0aiaxXVBcmhEPJHCOQLir1KVcTTxKZfZ/xXxp90uxXR
73l97wE064AGF9aVVpmn0zkFwZQLPwHwDPZrY9qKJnqY2KQh70YAShgb8l67XPCIyd3pSyMXYqRM
gbw3q15r2Csju/aTd8TQxL8MIKEp/QpOhvt5jCqa72ZOOzupx/HMa/YpoSTlWQ+vd/UhVcyzGKXB
eu4fj+b2BBHU1JnGb2a4vxlXL7pAjae3o0ceYwFbJ9LyfBdOVmjBzy7pWAGGa7QomffAwn4z99nC
ij3My4XKAdUahp4LpDwY/rYCiVFKBLNhUrtWz9RXabJn06AyE6rM51mY58lI3Myq7khQzLOkniCR
DlcfzD+c77oJf68SbzGjNKjRzRH3UElvdho5b1oRvG5Cgdtjr5lNT4wWZkTIOU7s/+L085bvoiBP
7urg/uzpnl94ic7ciEugFxoSDCbCGJNAeLo7QRdC+bDYJ4wYOx8S/5MNapXBDToOTRqCiQZxGzIy
+hiiW147bBUB1cR9G5vUfWftCdLZZ+JXcGswQfCZD/ASHprugPOrhWbgg3iFs+vems5KoR7Ro2oI
+4smflOysr2vvJdq7Cg0Y/xlRno9SoL0i9uDZrp1ZYgsXPswx+G9uikiygk1wCrfkXv466QaAEYV
nhSKNcd/8Kd9+r7qbsu6yaQQXY8pjsuLmaf2XcXE6gyrvH7MTUDtoRV8N/99wBemfQ7AahHxSa3Z
5grJvsRTW2+4OPyLMtuLo8rlcvvQi4U+75D5r/bs3piZIGsoPldjRpBa6dUnOhjgbwRICf0GQPCF
SZ2lwJlbErY3Sa7TbkFPO7GrnidOrCPgRILTtG2PIx4lVXyG+ea9Pxa1d3v3xHpp3NvQBWllbwGj
HBtleX8We3jmB3xnQwP+51T99LurPfa+6aaKN5oIwuwEI3db9F+yKJ5T1r6L3WlL3ldhbiwREabt
4ufGmDwGpqYHGcpcCdJo0u7Nc2pN4IEeazcBH7S+wVuTxY+lvVX60fX0sC0hIngcVsXFwleN8GYd
H8GTA7APgfT85rDjezr50iSM5+zT3cWoBQKibL0lWlWnRVnRiN4AtmqMCAUiv662zAzlSvifTZmv
Nq23ih3l2U9VdKnJCvsbyADfr/RpukdK4G1kW1EXOsB1CbqdnehZQxQeT3eLf8MiS6XQ73WmKNtf
RvaRsnbDJbJ/ePaOQimhQJS+qOkv4tFFBEk00hG8b4iiGjq/iAeQA9oN0qaiZeak4ZMW7bK4rK76
2+eONXjdfOX0BdNxMHqlIe6GFip/JxlqyLOorBQQMaM8rP2wT4Q2NPece8VJxW2RvqygYxbkCvLE
L7TB2Xkqceq8XwZ4eM7txMXLmML9PyeSyAVOGcbWRVpogMGnHJK3BTMHy9yYX7LM7L93Mf0fqz+I
qDOIwGci+XoxNMno8vDA0kHdV7NFd7xohFjXmKP5lanl9MU1XkVahHYUFbZQTSAPG+7dA0ujA/Q4
+tOiSagbmYHyIJaUDZ9o+kATD5k8cYyeVt7pIOS1ewncP0q+nmjNY+eOVoIQsxgDvIjmuhpRwl66
/eSXLTcF5Q3bOHD/vheagZopEFqALT0SshgYVTq0uC28bg4oMxDY8KFpHaziiyeZ9UHBqcmd1dUD
D+o7NEm+iCqHsLNzbyBsbSbJ1ZtVw1IPvCtpHZebfdAEgqXo7r6+gU3BDiu30UEVfdMUaMj9Cdi4
fl6Ty+qsJR69eutzKnISkmji4VtNCeOZBkoaqHVHKR1/UB245PjydyvvMF/CEXnPrgPqlRl1KZJr
4rN2e0nSGs3UGgmv0qeePrWOWZ253EjgGUdry+5c8MyJ4mTy/D1VumpXGlQcy09aFzS/ECEmam4H
62hoE6N70qVOETKmvPMJ1GU9UFKu1ZlvbeurUHc6Ac10f6I8e6AiRFVcMoHu6OyVUsK7Ntm59nNz
UTGMLbpNmxo2TVeTWoPcSXGbZFUtFod97pulAn3QQ+LKTy/hgiikm1USPYdNyIa+rzDwNVltwecq
pBo7KQ6COS1lneSAr/dxxidT8wN1x//rRzXEH06DQiAL4L+CDfMUDy9JLKcHyb7vo/CA+tMAomL/
PkLQ8klD4+McueO+Orukr+zFwU+2FJKWwgWcdSRhYwycNNxaxzbhRslk3cjBR5SpUPunZK4l3kPz
owmxZM+rSDSCJsJz2p6Ct6QDVolDDZ7KJpfMHU2VkqmAu0fXHDoMrOZcshRNtkZein9l02DGADv9
QltkXHRU2BCVt8nLwnNvtTFjRBeXzpavADuAEuWi8AejDlS+xFOd+n6HlKEZDKbIyU0bArhgD/VM
LXqqTZDPJuVxD3Xf7j/bWd4/qWuxqQ5gdreGLSqYUrltZA7qcBMDxVD8PKH9kTVe8gZk4BOiEJrb
KX/3qRyGMeZEQ5O1+i/8H3zu6nktuP/v5hj53gltW4AfR8xcr4qKnyFzlEHYsr/cMM2ghEd9I9V8
RFWC8t+Eeej9Pa1a5urd6oR5X9GD7PLBwPWnFetODU6depQXG+LmEgCj08E4CzqPkTzpkh7GdcHw
j6mKnS0W7LVhohCt3DxHPQlmYc+O4YmZdA3xT+TVPSn0i3hbYunM3PhiuaH+0TmHT1PRd/sHQKKr
WPWpjyRwbdxA2u2pqA9H0I9pwDumKkFQxlYePbsujXpt1Q39UtBO7N+a2ApFHE3CjlTzy+mzaxl7
h8MYxBywL09+GMYfmls7pKyyZamSepLxbYk+7peVfCXIeHn3LiLH79b0Kti6PWsPFm9KGzuz9o0s
1HYSpuldeBlLLTl0gnDDL2jIccZeGNV2gf+QWFr2sWOy0ljWk+KI89o2UQoNNtsJshyWTFGnppKc
WDvoovFgXODHADx0E3vZUYS1ixBoaeAaJOHI0TydKHoJRf0Bkx9V+m4RhnhfYpYrNH+HHV4LS1KE
mRtGOxYsm1Dd3w8UheupTByZTUWLp/GWgY/dbY4Qb6VoeI0lZpuvEXCYUgbhbZpPsDZ2Yg16NLG1
1H0muPPr4n3+972/IY8uF8no0YP1fsAucUPdgEn97vBSGdVawa/4kDGET+Njua6bVSmfU65bxxLW
uuTC766diQFkPfpQEoX0CzcP0CMUy967KXrd79DqsKmGO+nrUwV/tl3Z2Zj8TUDtb0owOAjlH3YD
IOl8avOK9oQEuLrEUXj7jlUZGVj/0TX6YTRqMzPQ1A9uDjUQdKUrdmtZb4KigcXNfIdg5DURQ8Da
LGL9OlbvjS09TYQQ4zjgCya/HgkNtfBBJlqPcnKWYZoPn0pBxf0YgQyTYMpd6gZEnYg4iseF4Zov
igw/ZZWcM1HO3/5MTXMiLrswMWU2rqL7RFi7JrJalQdQgi7nmP4XAIWk8DaVHIlJneTaHVxkq81D
7f/M7NxHvR+ET2k2r5orwb6h46zoQpxSySFS4CphP7fBFC/TpPyXMsTL4HvfwpmkQgtolSKVnLYl
mwIDYhJzSB67mVGVscjIYhRTZs9rJAGDXLzplFBkdJzMBQTg9dg/xX0vXG2OlKtLqyHpM4dVyMwL
nNgVa/Bd9P6usxPJzD1J16Lt/sYZLuXxmIMkxOX+wCjkXfF8MqthOD3jjPMMxpcniWmsWAgB539T
9SJzRU5k1SoCmZvQTxwGypC8FtB6gwwjvaB81lCquXVDKW/0Y/FFvHJfZq43dLgGvtCFoC56EYme
8JiXNKhNmKuQDiKYlw5b97v04meW4SevMg520mopkMsivPwZAj7iOHLAijlYvcB7arD6QOvNfbI6
yv1oARbzRluIaWh+ZL2QtyKoLm1wBoOhLqZ0UFeJI5PZcwGWvITcGJ/a0h8vVy56OIsdT3W3EQWg
SkXVlTHuTYgC3ZP/eyvlHE8K/yCMuKeZ4f4c0XgCtYW7n93DN0g2777dmXN4fiiphVY4yRnzOsfg
68elRck/dUH8iBs2u/PgXNNfeLWvSzk42YeXBpnYjyK5C8lW3Vvchbl7ZcemQJpZpokiLS3d7D+M
rIQcH4rE0wejpq93vof3of+WEpzVxUWpHaV0ARKSnDfXsejv3pfnfAyjxX1258OIIjtpU3dPHK8L
zoqyHQSGIL5Wxw+P1zt94nuTqBTvLK7hWZmIrt6gfIEAj7hjnkwB3+cbguMdvDG8PB70ossahyJ+
TkUl525XCPQDClYWzbB1AVicob2LAYFPtgtqEvWTsVU3dEiFCm5jgfBoDeNgIB2gcKt7om6lULOB
VgH7C/pPADOuhr72j44ekB3lpqDE/oidirAbnUUQqn8T0KKhJX2KeETbwzP+l2Pb7CCq9h8LhOH2
+hkbPUhfivhfXZrI926/6PN9fIpN1hSdCjXIvt9WYNGyTdlmBWOJC9vv81IjRawTtHNuUJAs3DSu
q2QmtGelE6815OR6/0Jxq5I+A42Qx5pqNemjgqr4NULIlUtJdXh0h25VX/uZLMqVYxg7AsskU6C/
1HQvIbx52wbkOXwhZJVKPLORfrAeMgsdadb82CjuQXNnLVt5QdUxK8wHx6dtvryMLe8B2DLMjPQe
z0ACm16DSfwOi8oRU4n0CTKtpq0vrIFvW6uOYWbu9nmQmpCNFQpqFipH060cXOYasvOaC88pGwZI
3EWtz+kQDxcjxseNKKx9XBVJGfL4McL6+amkAgjkOqnNaOcNGiGDqwfSAzMg82izMTHfnfXltfqT
7jKFXOjmpqJ/SF+PEZG7LVfSVjooEpI0Tx8Ueia8BAqyIlCIqShtJIp4C+5/pSmCRzJ+kBpnI48q
mg8I38iO0pTY0ZKkv9eoA9rAdkFSlWpwJq/vr1ZpmYJ/VR7f48Yprlu5JPaK8pUfH/Uyjd6OYkEf
sVKjYbsTleIfl0PRa261ZsJB4DzvuCejkNiysh5wuhS5gwtY8VFnfvDEXgnBzIP5Xu5YAlRTPUac
orDzXGT13KOoLs8cuK/D/HWp6MDvmVlTaRQCok2sk9QZYhrg7jKv4TxtjUBgYcv5O4xX0UktShik
h5pGT9kz8nYjmk7KsIWLHcs+y9UaXcyLoFL8eNd+S301SKm3fezyYi8WxcWmyrbT9fyVMzE4dW13
8bTpRmpzWxGivCQAF0gGeLfuAzpsvLSu6b7eaM6tyY1dNBwyrMum2YrA9DCrUojzQuASFuYMGXwJ
MRu0XXErmYJD3icb9UQBlgQGJQD/mo4Yt7SR35qCMO4oaL2hrCYLcCqfErw4/6tf9K7VQyojUIfo
4UNWTgHV5KK4feTZSTJ4MtcCuU3LZnHr8FYY9NIDag35qVeBMPNrnuXIsPbIRCOaxmMGgqLnOZDU
6LellDqJt6zHNt6Nlp+0n+XbVGd1uSYrL4T9g1ZNpCtj7EewFlAubVGmTYOaDouyrJOHkyyGy+qK
q42WtDgrWcE9EY7WXg2GY/WqG6dkeGTNHMLwwmMCi0dsBkx8cAsIflWVUQ1euXWDg7v6jC+GFHHb
KfveZsprHP2UTOqA6+ONw5f1Yt4/tAVvUVLVgsMcyhyfggpH9fZkobtBEcvYyHzGRj3AcJOX7Wm9
noKLjdLiO0k1i35Yka0yWbV7BTYtbqjtH+/8xbiMybwyM1/rqIYTC6QNp0haH1rLELnkaUpcy/ad
+yDwJBovoeljFLKTbgBuF9uqywIKxgSCiaUSkk7JJfKFrrnDdXzkKGaBglldyTzEqeoU26wlI/a8
WZOVccnWX4BkNjKCtx660VMlROlsvUgGbWgZMk4e+8fxnEvRNyt5y96Ddy1U3yL0te9vXBld+1mI
WLn0g01I/Lm5GUQ3LNcA20IcpJ25TqJZ+AV9e9k60zSNMo8LYBdZiaIY5K2cneoUHegGnWHma3R5
oGbTm4Htwtk/v2xGSiHvBO+IvpiUaUn8HfHoGWFR0F2AEzrIDV7HohN8ukH2ZV5SC+dW6581wYsC
MXsBFwXhEqODuccxVuzm5wnUVrju2i+2zSmP4aqIckZTYVXLrYhl77gttkdyF33d3iF5ToIOIhzP
/7Qxm1O6YE+402W2/HEdd4iR5OvNK2KEFNqEONQizty7qFp1GgGVPZC1DfA0gYgnoNAgnl4x6zOY
yVBEY5RP7dRJuWIJ+0Wbmg5gN0P8fgfLW/X4e+f6P03mPhtVSUvq7wRaR+V5UUkMoZZFpVM3Qd/8
tc3j3uX30YdjHZKfTwBs7WZBRcRgUK6uXfPWagNRiS9r5Xgpq9HB/gJ4lpD/2+4kioxGHVKdzyBn
CiFH0Yy38gB6F4UiAztMyGemwYSfmQwdL3xyYPbyn1YkudtLH/WCc5F1/8TFuIo3J7X5IH0H2Qu0
2hNXXxcP3pvkp6zGTyTwIHnUk984B+sgIaAnjP0496KDmVBEhfCk6ek5YUj3iO7+mHAO6o5UTgYe
UF2lx5936NIzmQjLABrNozN1DzxSEqiDMGoPZlmhKr+pu6qzVUjLHbmK2/nMCb8v8hwDCNg2s7oS
1tCPjnai/Z+GGzrbns2i2P7A6CspvZqwEJRNMgQgY49IMSUvj4T46W2LMXHuud0OrxFMtpL/E7QY
QyuwnZWRltbO+OJAzxTWjUmfCyw41jTqPYsCXEIIVQB7RkxIYxD4GMzXNV8CU9dDwjVb523a9QX3
NMwWt/OWOrGnLTSaygU3HLMQu74eygh4Hjxc+Y/25e/Xzd8EuNdrJ3VaeX0/Lx5PQg5lYkRhUC5G
oy/dIybUOV+BfGhgNEBRCNu33qj03kATXwLLPsio0N4BkKL1XsqcGw6Zz1wfWT1s521rMfmGyu0h
7G+UrcmhlXOaL5KQu286A5nKpuADleEpsRJU3BNc9lhJWYNvCbqOdGb1PqRWHzJTdYnWFrZYOVZd
SAFt/TtIFNunZ1icWcwh9j1kVz1OI9Q5BtULkXDNumG+PoHanAxzlRDmNFOj5XF9FvZA6FIj1GVh
YjC7raya6PGQUZI7SePGtTwsppYVHRu3QKot+GlqeUi1+q5GH7oaxzvbW1mcB7EgGmQ=
`protect end_protected
