-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vIXafIJaseZjOq8XfhGGnzmM1SGBUYueOHMpkkRphFhElJidJC9fJI2mewkeQhTwW1Y7rsMJYeg/
lYHCl1kk7e6lA7q/cbGyeJtH9Vk2uPZy41labaeNdj9oaucuuqFEIzjDF81XB/5UuHQOzoXqcJkh
1PXBhTJAgQUBv1MaUYmXD5/XskRkmHG+Kf1l3rAfcFWkUp/BbVng4MLIJrZbu263AZhCrjQ4VHPr
OAbGGU+KNl/R3N44mmn0VnUDIQMlXVst1QM0YakKf8RA7kOyz83sz34fTbyc/fP79fjt6GIM5R/4
RqvNa0KTaN25LZPkgo86slt2HpQAxy6eHe3tpA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49216)
`protect data_block
Yzu40wEXmnVFqEwruZigXevOGE8uUsFB7AcipiSvwf9t25ULV/CN7siIEnGRyWF0kLCZ4cbrbGNf
O1AWzI28oDu8kz+6OdU4yeiEqM4v2KH7gIDObAFNr86GaMJaofmAIW7x4Nl4WI830wTRRUQYr3wp
V29MidOTlPF7iwkVguhzYhTvD7nVCSWk1tYFdJjHIeaxxIuYVlGVBL4csoX9y1h4CmcGl1+n3aDV
JqljvNQ0Ft2o8UkCxO44oiBgCyJodb0GP4Wav1uBzebmcrYy0x5MxqZuG04bnW0YW7fRJmF9clow
P1CyIfsmOCi7u7FnHCpFWRXcsLkXzu4rb81jyx7G9nlCsz5Oz+6rVTOW8XY+j60haR9IqyhiQiwG
lDJayqZnqi4BVe02ePo7QzWOdH5D0+hkBQU5ewiq6lzoyir+KXVctwMFr11cygMhBanQHIHSZnJ1
qbcr+Nu+mOJnX/5Tkaorux402jsCAs7qlEYFTBuPla+TX8vWKfqaKeySuzFyU6IJ2Hv9uww5yg4K
SN+16OhpLm8Jk2SpqJKWTCde2rvNi5NVSdLB9AGT1GEv/yNs/lAmMdablPNrOmT8CwnYWUebhy7D
eOREHb2/7xCucMQnOHTt1AWkTk9iR7f5Vwtv4/MpaPerk+FAN5y+MBX6hWswY6IzoNNYW/Lw9UaM
BYWV34x9vTBrzU8GPnVBngBFzwGihPsCPneLdmoMZsX828w0dk+zxXFl3XFhJDmjPFp/P6Vn+V7h
jhrtkrlhWr+IpEt7RokFgBez9twSv503QPb5Pw9R2iPj1XH3Qxz6lXPDTm8As9vYdIP/3dc2jIQ5
zriveazyl2XQf+QWDGfnkywxqS9enhacSbgbKZ/Uta+MsA1EuUoT5PEePnK86l4di1sbY/7IRQhv
+LZnswZKJE67Fz/cTuoLsDVGGaz3i3GnBZXYiN6eG1h8v4hdgXAIQ1kUO4zw3ikU7P7thSzY1QDD
RVk/QSgCJ7qIi6JR0LlZAJXAwyB5PHkAi9ULxWq7nviDi+UkQBpqCUFCRmhcbKiabIRFb1a3KrEg
SVg7oirv2ZgFt9unNkkZMwn3n5moj4b+gKR+g7KFpHCS/QgrlogYrWO0fE/CL5WopHcWtUwFosEc
VY0G58vw1KRCImxBBLVONEEb3rcUcpLR3OX75McqQt0T/bun4HueAcVNwThugNEf2GbeVknmgedI
IyUcEHHHKFNojf1ZLwkGl1Ho8P0Z+/c7j04w9B9PxV604lDo+GTDcNaZFZlaQtevC2BhEQVzaHJG
sIy8lDRvxi5Dvtr9zRBXao5SlDbQY0d3QmyYwGdbPIIYlwNRJZSfGaY/YKWve+qHjzzWggx3p5VA
ExOTr9yHYjcq1mmSp2FniPJS3WKY31HqzcaIN33DUU4CqEMfp9WeU8KS/NOP2pRczdn/TQvBizpj
FoMwA5+bY6tua36ueqleQSOV0YAS0CSWyGkc2rrs3Jj46JL/Uril+8GtsyJd6x3e0FqWhwa96O45
n1j4jhlIIzjKd789RZ0SVTGMMPk2G2+evVDQnfw0yX4y2DnmH5EgZEjFfbRADRxXGnSMelHH1DyT
VGBvbBHcGMVeuV7ShOuLDO4X5iExqx/PPmQ0Y/rChHry+xODDQuC3rCk3JYvZMZQS4ucuBbg1DPz
j+qi5pvdwvfdiBXRdW82cnWg70/fxYvzeMo9pMoAjx976VOphzFKLQM44uyUaCxpu/WWgB0YIWIM
cjeV58GbrKpl6ydgzXkrOPsSEhBu/rakBPdcXCHg5V/Rl4gSdVg62W+OUDz/5j79JJCjASlOdjVJ
LShl20pXOsftakMPQqSM41f08HrB4YKiXAdfo/+WyOpcmHH3JY9LrBV4Cpv8IPQ/jodSJCr/rSs7
HDc1Rxe19nWhjMJqc9TV/zOnc8tHkA5yYKAy3PJjKSvRQaYzVMaHJPUrQgtW3eVAvw31gXiXENI0
EWuVMxEiNC1rHY5Mrc6YVEHNW1V8+LUHGrcKraF0CokUkYslSA95l/HH3/DvFRoq4dMCNYx23Edm
UBhq7s/G9ot0VBst033kvNNjgXRyqh3/6lATtiPnGx7IEiVn0PSF9J6UVWqrJdn4Cx6N5/ccAl+s
gb/lcirGaUHA1+QmqzgmcHFGoZRDMcFftIzXe2rpXqPBornEykyo536mXWov+nIfdN5E71IH2EZA
9u69DSe6/FL15G14YW7LSddo5NlCw5pTvV0T0vrSDLnXpX/sV6ba093lTz68etNlEcqH3+lMJB9v
u3C8jXyMgV5sa/hP7Honf7IKf7eZPBNTbQkAbP0J7sVMSyLdDV1ltDs9xdWmcfcRnPOecVJuGqEo
qQgvPmx5sfoI5sSPFafp5DS2J5UPKHNTqWxsk8EFCBnyYFdoHVIHM/khSXbDkYLRkMcCzYXNxvMO
siR3kIIzaLkFWWNrQ4ocDfznAgAVtGq1/bwb2t7zWWmnq6jz3NEgMDQtddU7HLAwqEh97JX8Rnty
wGiKGMtr3FBeD3m8XTkcgmR/BqM1+ca0ZeMZ7CxcF7AssTmRnZBrAu7zUk/hIi8nZ8V1/Dz6IM87
5t4nsLS2C9w+HRw4AXLpYztDAM/pYpu1Q9LXsLnJLWoWk01wniLglHxMbYjHcRbdKl18F7WwsWsn
eEQ3Iesx76CmbQcECdfNQzCNxSxMPf4i7ET0wvzTjjhMbDBA06czxUjuUgRNjk5iAw8YxSnIk1n4
+VxBBY63TWTYGRs8IVMYCD9+yaybpxqHkFSlWYKYNbgTHJ4+kB0bXyo71PLJg5qQ556qCJgejOKc
R60rjQgSP3G5trKSJOR5UVOG4pGLQAAosR5/qQZrheyR0Z3r787QRDUiA9RseD0KEYxhm+PT6bqB
ajLVUINKt85H+C+K0x8RrhzD1gD6bAORxoCOkP17SxWX97aN/3pHvCfLH6rZK5QvjwusGRwiAifn
Mr8+LgUFvAAx7eH0B3Kiueu5esh1QgnBmvWQnYVnEZX98ivBfayryrliw2vxTgQrUvuoj3IwmLQY
MocivyBXoWhYP1Pys+w+g6MVXk4v4Qmfz/XgCMIWGu/3hD86tIGczkuAqRcJYvG/l1AURGBH8W0Q
snj3Zq3atB+4JOAXgM+RR2H3u+8aUBs/VS1/8HFDmZj8U2nNKu0chXtX4aazdoX4Ns+nEsq3j9ER
qviC77kdOOmeajv0dPwpm6w7lUBGzhxPWislDwP19DGVElaeW3nlkQ9INtnlcuC1WAN/FOTKPJEL
YJv+io1e8gsBXBQQYowxIslY4LUkdNXLI4fzbLdz9j2e/pBvGf/BOfT74xKL05huubnD68ys15Zn
hhoGaxxWMhgj/bzRP1CT+4G7kmQHjGeqZbZ65XDlNzNeNCwuinTwl40NPS0T8cgg2k07xgQE48gp
QO3Jk0FmPlJ4e11LueBeQzTLftBvFxew25yVSsN04hdL+BKzl3hAswcASzTIRNI7jgLnN/anHZZp
7hT5Cq1rFqz19639kow8rWjzQZ5tIVQmPbTN2z7L8eVYsi8DCoMJ9UvUd+OqTtbC5JOO+j4cwrUq
Uof2fYuQyxXOjKNmWDux2Ygl+UvP8QSs5BFhsP3WVaK8q9MPsaq8mMWC1BLgQlPPbWiw80PlOYey
vZvMV6D7s3jv8vSl9qjRZ2sfb0unHIJ77w0ErkbAw/RnzVg3aZO4sLTXWQHZHGzMjWMbTysbdOjp
qJZMp0HK65VBVR5ZpaH6jUcReBunG27Iy5mJOukiruc1ub+R3PNB8wLnB7r6lyAyZrna6MxMcLfs
mVif+KEmuFURrx3/DGUCDlceMdXwAyDO7JezrO0pxWOtXJ3Evu1LXDauUWlh9YLutQA2mXe2Goaw
ptf12coyXx4RE3swLhkQ++FU2o+G7M2uL/96W43TSBwZhpyAt7Xt5urCcJqyKiUsNzKVuYh9jLZi
VZ9oPaor+C08tCeGpelxChoEe02OWSvf40VqouZ5Anb5+z2xxo2/otf2CzyWcPyxLFEO6zCkqu8i
t8enoGIEktwgsScsc1AYxJzVFOFzFAcgrmEz6F2b751wParxeBYyVPWBJapMpwNrGZeq/GQtNQlW
Zh/dAGpeZPSksd3mwQ9C3KTSOlkJCMyCB6+jaEVz/mZY2fqpNjlf0dYq5u+CncJrbsXChp6V0wbC
6UZPNDqBLELT3YCvlcozDlkHEVdqjWHnTCvZFeqwsE6oQnMbIQvuHV1TOeGjoeuj18I88KvSh3HR
n76qniQuEE3PKv+42pKNCmND4dJVG+liwMo9/P8ZVL4EJMRVZ/gOINI/yZyjjR1WfRvzrjWueyil
8Ge/tZk6pxjGSV+elXhcJbuyIpXJ8Fd1tg/IFqw1ZuWBb+DzV7I08VlExjOXtO5xAjLkx2X6NCga
C+4YUqEf4L4w1gipRhf9jl7DGJysF2fT5BIEQvJ0xE8bnbkl/rhjU4EFvlxbMZknNdwHn6uYDkrb
ejApyuNCVJbUKl8Wi4+4eeQDWV+hM8nnBgboPK4AQIFKkxnxGvwIudHJtNJgpsXuDY2UcEjXVtuG
IW3Ddb45Hh515R4d0FqnJe6j6izPp658IJcYEHnMEEWspIrAAZrL47SwhSsHG7V+/T+suRwxcy0b
jhGJxSBccd0oefCWka8Ri28w2vMlKu1duBo0+B7q/gw9ZVyylGCUB5bb+Z1xGpso+vtCiDxcs4v8
tU6H8TZ0j/HJM4x+hkLwxIXcDhPq6st4TrOa4LVUIKMLBmpwTwHluZAhWKADt2KFPkBynRHclUoy
fZi3sq0q/Na/19MvN+qx2JiC0/lw9R4auuGMXL6kw6irWfq9VnMj9uFQkE4GPoLqAOVtFD+JFfIc
zsqNQcmlq7Ep7AWQWl2aX5fqcmO8BUy0+A6sHjbxkKYN554mOrgDY8MUR4da1Ym9djyK7qLswiK8
jcbhuIeJrn/aMNQG5AlPbUe5w28kRRsmvpoBDkVNIEY3tt0RFivUVmwmdoIFgWcT1RMHENEMZBED
ex5yqdIrJiIF0WWyGpOSSKYHDSXaPImwm85RyBVmM6NED1wVuec1++lzFxPRDkuxFg4DYX/5pvuT
Sp+2QZRE7cNNdeyBWnFkTQwN1HKazOaeLYFlXrqu4zImeSo2BXrly/lofpqLawaG1+6NvTew3AYk
nC3K41gfy0hoeJvuwuY94Z9F4V4ikmhHLXJluFI2gP+HyHFi27gexj44pzLt2KNSYyuZq+r+UTpc
iL0mWxb/8k0mPYhafPdk6WTanmevOO1soeXQD7bCfQyUisv9UR3G7OiC/AhE6OefWmYrteZtsCnk
Z/hzYud5D0CpTt3T6jdymYXATrZ6MUULICi4SWQl0MCj83w7pGYzNjZHaEyHBXePwkyRL6Q4tjq2
E/c2yb+RcGrEL3Xv5+aTgv0aQlICtRSgn7VK5y0dSLRbZN/BDNRr+LuXw64JEVYn9sEJ4cGd5hXc
SIHvTp6XTRU77AHvCCfOJxiKb2//ANmR9yYoikfa9OfjhPDpZlcLqngLSkWFXTFIGigaeuEJj+sA
JEC6FAxswvmMBR5OKqusU3HltzDQqEhBZRKcveLqcM4toELEbdF+YO92rQLcpm77ojwiUAVfBFLZ
pmiD7iPQ84LJvrxo4KK6t7jg4FuKLkXNH7j6yLspWRvTHvAt2zXEdD9DMC8JRbdvddV9gt396IZN
GiIaA9wIjY2zHmRntEGWtGf5yw2mSFadApgHjGBvbQ7UA0KsbdDJKVX2BWFcaGNztkxArqyuEdJf
h/wxbHaHjWn4iKqErW9Qk4BEJRwUS5mwg7xNQzG+oXcMsDLmGFwN7MN3E9ddY4siXXxPc6rn5yVb
iCEHX2m0I8jSFdoNpt9YNkT5Ko9bbt7S3bhJ+eoZVwyPOWcRvU6eTCi3Olo0pc2x6aUQ6JvcbZ73
rgY6pjk69q45LFEP31AikHXi9ekyCYrR9A+Kg4ta93wC5p+dylQWjElHtBh2M1pINIW1031EPio6
Dw3OcM5wualcUkkiYLGR1zp2NHB9E4Bmtjud0mX+eJyrFSEG2ePN89IbVeHNzd25wiX2/aYKnUFl
LtKlgBOWDANjKVsyMGIOjLJSv37+sG9ixfP98/x1uIo66GbnF9kBS/RAKHqCZ9jPj2BA/UyyEqrU
fW2SQWw5cgzaIjm0qZ4LIFtNBLcrwf1bQEGT4TLs6OE0deH8cMk+c7urx7f8J42a76Ca+UkwN/cp
FuqPqPVmyYxI1L/p+4S5VHq+hS4OhvVdiHjFAxh/63AN4Y3CB3GROYpZwHrNN4alkaN7ONQiMaWn
wRE2KQcgKI2gIgXRSdKe7IZp8Pa1JdEnB+K8Je+h5rc4e/HVq/HsQm/fQmuHTaC6/zIZ5xSHg0BL
njujdGc52KDKS/KqLMdeZ2KtkYERmg15WlFrf70KWn9lYo8U+HRXPdtpyX69Je0IOb9uXo1Gtxx5
153aRREYxp5n+TTF3xKjffxCBTi/sgTgOlYjJOVJsAE6b7PDAZUKYfMPLYK0i0LrFVna98lMZglL
NGAyYLtc9OGtHUS2H6+YL2Vp+ZTIKhLZm7r+5t0oFzQvZaUbXIiDnTRIq+H+2f6J5/eGq6uNsCVJ
2RPX4olj4jQzDn99DeE+bP2bQZx3MBgK0sJJ9F5XZfMueLNWeVaIdRlLkgHH8mWMIn37ZCvwg3Aq
jUDp8KjH92URlpHTun9mkOAlR/N+yxzH7C8guMaQ+beHkQojf+qMpF3L/2Xvxwdcn6/C9gWXNjwf
PXuBnoIC7peawebI8k9cOyfYI2tbQfw++CBarnFLbQ7XyWqyK9FpMxpOIGeCzAD4u+gVfICHtbhY
1hIBTlPftK9/pB+ZZwkONezxDySRr0nsqCuYHiqUXQtfiXiW05qWIOS0ukUHWxaL+aFxvmChKUfg
oTnVN06mQZKiMJnfYqnfa+E6Ah1OTLw4ZmA+t6dMgCEkyPJ0gT7IC60bmUNw4YGR8bQfJJf3rQmu
LRL0/lNL6L3rDCamD6ArfvXIhYAe5hrtm23sqGsrTK/syFfEy3mcc0eN0C11FkhVpGVGE3sXZ7Cu
wjjR4H2GdDxC2A0BG+Le2qhQetwuuhyV1HudQ9voiqybGgeZiVPGy0oQ9mqIOdmnF94k7LwZ/7ua
3F71AOZBFlSyEUZHVmS48F7JDRL0W33GnlywIokeUcTpct8jFtXWOlGxelRm6bA562ZEhizdp+JU
bvmSnsNTbi9qV+uZWYsU8liTqWf/4zAIcuPoyo98vn/eMANJbOvTgky1e/9qlF0rbZH4vMNY/XAU
ft4UAOdprcYzz6k3FMfPIBjcADtiJTQ5YShTG0ODdLs1Bm8GlXPRayRuDSgz8U/fOjAwRYmlqEKx
hcWq7/m3XCMl5C6s6pUhJ00QIRpaVFL7o8b+d1zIvRSOCspaf0JcN/Qvvksd8hi4wTkbAj5LjlJy
40ubi5HcGRPxzqEmFJR926HpeGZ09HpeBYIpPT9jhGPbw1FBr7HlnStFAJhRM/LcCoXHb8+MyaZJ
Uwq4LVeqj3K1QnijWbSltg7x955BOkqzfFYgbCHunpoxjAV1mSVNbXPkiqJEFvqadgfX5srEs1WR
EjYybrpPqNOfctNZlQ+eqxXaze7+JONnU0ilBUj028gPcAOkFPaQvJ9BDl2uZGs0C9Q1iLnYRt3p
bq119S7lAYs6olTzyPciBAln9lj0h1ueKJ4oVdoYNv4E6bVX7j/bghBsZ8Opeo0uVi52Heav3QIF
7djASLi/rPzZBONnJaQcP9dXXsDW2nFwUTl5n6EziINpCSjGZ9xDbpB6syyRg/PQl8LUhSDParFr
/PeP8nFHIC9NXGCH0wqHudhmONyrfeGQHI0EuFEo+4EKDUdlMr2sm+ir5hHG4gCmizoEU7b3Pvbh
mLFQIiiXBI+joUa/83QIGBfWIFQr7aOe3vukNtxpUDnX3aQJcl0k13YwzkLxDejlRXHZA+C5gj19
ZxePu9G0XualUpBkkPyGhg7N3l4ogDwoJZXGtypbFIbcwAJTUK0hujeegYmCbaZ4LqFPAgCtttHH
x/OjWJL3o1/xlfib6Ss2Pe67sqTs99hdzVTq+zFZwz/giV+4QikGxebGddZgooGVmdVPCsVioYoC
GnRVIpIYx7fZvtsUoff+jb/eIf/BLef4fMNaGkK9dAFAZExN9TRxQnZRgl8S8r/fiXICFZBJk2dk
xMrv+WQqasyvylyDnHyyIrCteiJpgwVughq8H/yPnhWwGJgi033/ZdygxUob0ukXrfvSxyESpNJH
P4bh4/stm+9Bq7WoPedgQIfb1Jsyq3T1GPHqVizAqslmLYrt8LTNUEMW2kacqBJ0bbVakstEImYC
VcWtGQCDcGxTf32Z6wXYPgBEqtXjM/g+tnTUMHKO/uJ6H/sL3XB1BdDm2vizMToCVj6OPZ4FpIlT
+CDoplYrxoXYQkSn0nfSx3lQefQoTaLDVa52GICNBT+t34C+o24vDhppsiMg0xLv/MxLWMmWccjd
ZqixPeB/LpEkiUofOrwQl82IT8B4L6ojqZAhKnWKfg5lmb7+RN6rTVMycotRJJwMpKCViHOH/Hhz
iAvZ3RsyXS5Q9asezcsXQ9ZrDKKuzZWG9XeWvoZESeQzRWoTYVDxbfLAvKlcmYqPvGWSDQzZto1e
kRFI/SxwWPZYEOK+M7gKZUGFGLAfzBZKnkM6flSdd5OhCAD0KMAwmpin2dzV7mHrRj+FViJakZMQ
nv5623fsOA8ibjApUW48fNBo1pFWK//F+fMV139aSRwkuT30cJibkmjfe65HW0GTrY530eiHy7gQ
GsxiiQQMIH/somo1ZH90xd9eYZjtbADP7Ai7IX41bCsZyBCyCqcJgqvXGEfMOce+e7WrGBUK6OhA
w1IFtYbLbokFfXZtYZqC8ueo9xESaPLUCGrk6hWEq4HAVlQQI2O2/km298IhOhKD2Kqs6HeeiGMd
/x+z9yKpfqMuWbw1JkeK51QuXJdqwFaO4pOPin4jX4ZL/LSrdIUl3UEQvnhTQcBZj/L4EVer3E5H
P7knjVjOxUMbc0hvOVFq1Nyc6CzHoqGjaSz/lcsgrL2owSoBllZc8SgkdJpwx6gnBZ1FUGLqiI54
INr7PiPtOWLwcp6nDQSM8Qbhr0HQCSkdRRDTYUPqMbWLfLyV/owonsC/EWVd/B+eHecILkGTzbm+
kyXdgI6wKU1PvlHPUepknBAa9ja7++SPA77BpSwlq2+v3CFc4zIqIhyOJ1s5KDuZ/DkfLW7p1MgE
l57KvytzBCJxGH/pbB2TJ8znH+NkD/6oSacEE6kxL/cI0hQ3XAo/PaGCZfxd8Py7aSFfM+ZBCIQr
Ci/cnyYpEpqnHn53FVvk7bV8OsKt6CdPcfATsovw23eKZfbdKdPVLNw2Bnl94STEH8pIMIt6cPRd
XxKOiFMMVZAn9avew3VUaWByDf+0VjYrrGefCJ0qL9rlztLYRfBQ76/ue3uk04VpWo0IM6rCIXxH
ivglgXVBOJ4XjCJTPSPKDhbiyOlpNXVcLoexc5Jy+54FJEz6PucUa32a7mG4wrNnvf/f5CIv9gUK
KdwMbYYznCJjdhWvCy8lNWeChYevYWO97PeJNWjg9h1eowjD36rO8Pg9UnRKL+SWr/4LooJTHaeo
ImJLzwXk3gd2gVE7d7NvwRde+K4CQ5zQ95jAE9EUc1d1+Lpmr5J0Kpmqy7FB/oYbmDGZdaVZkDFP
Qy/UVnNsXOYdmF+NTWEl+pGmkERq9NWY2ydApyhVGqzSze/EM7Hiq8EbvSPf4wOywYm6q4teKLQB
Jr3oS6ZWVqnGSCBtQv0cENh9lW6DfX+Y8rInF8aOk57fibpZnIfRQxS5poxLEPz5dL3Oay3G/0TX
1DgMh3Y2w6DxYOXvCImO5ZuuHBB9UgcW44lLL11ORuVMeMHeASgT/k6LF+V8/mdoWs1Ek/5EZsem
koRRj2flCn76e+b28FyjlaZ4zZFPVae901f44AxHkFmkI4tFV7hdGgIu6nIQeuLtuPUCDbPRYmJd
WAUI5LSSw2WgnyFO2ilhZ+tMpjnta8tqJJBAXunFVG09QygwW1rNbbHDoraqbg4YqFCh60WWq5yM
9aFcRTB9bv3J/4B99rck6PDepeaZwihe07WOwmH9mX52xi6YoC/LS7BOo49d/NycUdhb/2EuP2zA
0+6RIszusC5EFYEbc9KfG3H02UNH0AIgbgAiIBSRk3el4ooNkUppZsnJYgKN/jO8JHbp+CyG9A2f
xXpajHs6uS074i/KpLEo8iM73XsJ+iSntoauAfBlUeCPsL6EdaIGjY0EGye3S1aA5TBjDwM+0SVR
F1QKTYoJQMgkA48K8xmnHAaES2o1YMZpGbrCSX59G7gExINaz5QCE5eYkmD/mRn7hkqcIJz0dIpe
99hyj2homCWnz3z6ldU3Htcl3w4hyHdHoTn2zAE3IMzCCx1up1nTYzjxoHXQHdilogm1HLxtttHE
rFL9rHarAZ/SrvSm0dB6sk5xgVgzP4vyKFHxTKVTHpTQKkLTSWTILcH4kP6X0NxZq3uvaXxH44pm
7R+/uaikQvxAKfN7nMEw56HP3FphipndyxiX2+b8Duw/YfAIenwYQE8c03fXXsMIkw/GzMAACRlu
p95xM6iHLOGXWBD8aEZLLKpuSkdLFmdti1ZxF0V7QTxqqY5wLuSlh9AiZAcY9V2C4Px8m+fFvpVm
xR5hNs4ZRQkWhRkQkS24y3IV47I7WddH/4Fu27krbclgfTbSG/fRTuTiL2XQvGW4RYeT2tVN0vwE
Fe+RLQuAuso1Paswp0Ot0ZtvH/w+eA4XN7PCR+cCOUVLd1ZqLN0BuntyMFbA+tHHqgLhYKC9TTeF
k2uKm+NmaEMtQ5aSmG2lsPNR88HjawWRkMnsDeILjfLGIcwaZPjH3bpnMzT+pG7yDdQeuA2BYmAK
+ahrsjwzJpGUXHyMi+9Bm/NniANYLzaNT2i7xeYbSXC/Wm8FU0yg8lZb80M65nTN1N27GzbnoMzM
YdLiXSyQJUmipy29Zy6LgDmK0ou7KEeWal1GSHy9/wn+Lw0gmWRxSb1zuD64rR64yP6MDp8Lcya3
U0jI8cC6cYstBBCAYEtD3Y+LK5wtw7uu7R+pGtfG09HJw+aPL0StLnFH0x63bhNdPtZ8ZIyVLbH4
JBO7vtAES0enFkOm2ZwJ7CQ99QeNaA3XXOGP22Tlj3zyXKopYuHrkG9OGHsc2/9yiNJWHmpEhLM7
ZOn7URP6C1//BcPkuT2lWkRStSA0+mky3b6mZUnPjltmmFOduTUyEp4a3o7did94rHluBhVI/XWQ
zJ7mw3fZhLu5ZZU0LzfHiDFrnjZPLEhLab0WxyQyrvJE27s9ZHJQ/6P1mtD81dXEChQOac+spsWU
Gqib1qGpVqkWeJDvVQyoxS7kfQk5cXldqgRUc3DR+z4snnqOHjzhDGZTP5dijufKzaaXmc9F5PPl
gzbeQLIxQHupKQUksQomzYcq1BUGUeD8eFrFJrKPgGvD7sJMeEhUIRWZm3O5ozeE1noEfBon6fXH
X00VxqJn44Z0t28ctznHsa3fbeA8H/XnYuYuIdwdvpy3b3tVF43CmCLD/DWiqrXFeAmlWpcjYOAs
FM3M2HiPMhEiY+D5Fk26T50Q36ICbN4l/yQcOuoJgGtR2Uhhq/KeRRjlrdtXoP+hZEjlCXLJ0enB
pBO7RoiHCJbcB9SmXeyD+R93Ijw7mwt54PKo3bS+JTe3T3GwkVWoUSVFZe8Ec2o3ucKDvY2jiKKL
0dy+tJNZ6UZ2xvvvAd2kJJtbJX6Tm2gNn+jClSgeEgM09zeqIjou2bkvk8pwd9IzR8Z2HvG0n0iW
Tf/KrVSH6ZjzNhzoQbcKobJn+y212vNz/zaQ9M4Nsobnvwqk76clmK1aNZNhBU6HDWszM4Ppvc4o
nlp6slOLrTU8/QL7j8lJleD78uXfa74e9X/sc9rqPyr9PTDJb4xI2w54Xt1HRVWApGTlbnocWFqm
oBv/OlgLtzmL8AGzxiL+7KlV9r8gVg/D7FZaiXkUba4V6L2evimK+wWVz3Ga8ngZ6c7pDiYGH74V
3kzP+f0h73f/H6v8rvmvMnsoeeMKfh4ohN7rmmfRqELhK4cbd6hPtS77ZEHAyLULwIbPYCclL3Mv
fq8JbwlMCfZ9fNj1ngPmUN2H/3cAPMROWQXxPTNgIeOYRZg/Pp5zobys6ZA0KMhXRvp77Stw+RBn
IDvxoVZn4eAYxk8ZtVb4l+D4WSMM3BCmTrCwoFJwXuZFsOadAIj/VQeF3kuW9kDdfB+xhue7dqLl
4OF4tuJzpM/i+MxYjlzj3tM6hhgX/+bdIud0fA4orMVcVhR4MY5S3+IWoS68S7EcftE8Dkhyv+KP
OhaibYBh8kUTGraoc/x3KA33sBUXep+mNogr4NZcrC8YhWJXxYwEYuj7xQUdH7klg662KUXLBuMB
nSB+gs0kIN67n+RFOogw7uv5bU2Juet5ofJ4ZqVKy1lyzDAdE7sa44TseFWa/iRA2sEDhTmpdWtu
XQhbD5pEIKMMifHM6EfJNUxZZ5eMxNpwtG/LB1IEkcxnBU2H1qBr24cRJfG6yvhvkz1ZuUXNjfJg
zvTB/RJmWSsvmdhNkAs+NeXyJYeUm4VrVPk9tfQgvZY4fdCEY8b+auSPgDgB11QqyhdGSlBqkLM9
rPRQBcOV7iUMGcIgAvBDYfNNS1vnYn0ehGEslK0gOO/uMI4Zeq07a/+IUoO5ux/uDOFZ5RRaV0t3
PBv0aXIcpWus0e+KImgBIy4K+GCMzFWJiWXbTCvlx+m213nie7PbWnuAdTE7eGrAb47zI8QmTnXR
LoXfH81Bb4msbqDATYHaesfDjda/8U1sUgSssM9UWUEsH6+trJr8i3D2ZXmChlloeCmwlNXc1bsh
OHqJGEm2HUhUCMYA9M54nsdNeD4YKiTvAZkYkiophZ9i+xy7RgR5og9M8W9vxHtkzYjzDiWIgWZV
iuCr2yDG/C69aQKvfRGZdqw5RpXlvaFEIJnqybzj7QCoBKT+AgBOJbP+o4DAcnSHZOAIo8sHLp4H
aRL5B2UOPmim48ZsQDBU5/rSg/YYj3zm6B5MpU8StORIhdxNF/eaCIRmYZcweSlGWZbUKNcaWh64
StwjAOK2d15MTc0MY18/04cMRqtQLteB2lE7+1faHgYKxJ+djMDgj3wpUOeyM8FmzJFjgFAyBJBr
NlXczs63001Egj9yTEh+FrxjV++PQRZ4aVYOxIg42Jq5l7fEHiYE4Vbuv1QtqJvVltwmIhqTwhoI
DOKbT4AUj9CzkAbyJFrFjDp3y4XKO/KObpP16VneZ3Pdj6USDrSrxvaCk782GNXg3sdTZIe51e+l
D5H+U75Fq7hpB/EVH6GA8ASdeXOcnqn3BQlsrPaDR5Q5SXxKpQWD2GlHlGZImeCyieKA0Rp7Hdqx
QvkJWFEDeQuUjhb1RKOPCFyrOBooIrP1eJzVCwEWuDt6xMNP6TYdY0cwxvbPUe4+Jf/zsPOZvtnh
NKEhiFqOviAZr2Y+4Is9z67mdLMZ5ayMQge5X3X3EvVQe37qGUO7zZnXNlSWYCJmtN7wpl7+Cfux
cyuIZ4UuNteTlHsy4C40N1oCHppU6ZLeRyPZe0S45U7TF9ZYwZfH/lCFHGTW1EZhdla2PEqH+Vya
2o3PzovZtbIOKw2fPIq64+9VaGDnKfIhJcNXh5zBJhSKyL6URdzh9Qvh8Ccu8ivxZEfaXK4PCDLX
usuoz5fg+eFZHBUDqiwR+Lnb1s5cRxqspIJzC8cY5an5QBmAFp3xkyKVb+QLDB0U5BQK6V5f4m0X
uh38VktqAVOq0SbK1vFYdOLET7su9eZobvHmSWnwzPUsMq1qdlSzuhkpYiiMhT/eJULF5XFLKutg
F+JuPcw8S6kVdIYkHZVTqZh/kaI+3Esip5R0PLn9XpicxErd+kvlvPamTO13XTrrUWTszMu4ql35
YoGu9Jf/h7yE7rNf8fCt3I6cwmfG0R8yW5KXdhQgawD7/CtN3b4aJ9NBmqbKMhGD9dmyQp7tvwW1
FRiD5Nt0MKFl8WHweV2E6Aa7O8GpE5jwRBlquSd9ss2B3GEyTCvE7TGsgC8/tKqhzSGG59udkaCP
lchaBrjugFmGsfs2W+KBqrmXfV+8Dfa5Wb3lbdTl2U8j8HHNiOwuidJk/hUxXtwIoGKPCZsLbWJn
cRfc4jwT9w9PoE58QfditHn1YcaRvNAJd1HUS1cLpvywjgCW/OY2FbxnFlGRih5mpa9mqo5LEgYm
GyQgoId4nv4LAA4tL4vot4LyKnPOvD9ul0gREMgq8FoUDA+y4cIiYn+fZyHYVKmRG6HQMM836est
z0Z+n0mmIRKxKAImGSy+Zfd/4u7fiHMXjZiW0XCo/9FWdsdOcDe4rMLAZRJQmtSjwZVin3w+u1rY
MP4o8IA+5ZzrZkC+owpGLBVuuu74VFAJ92NS3hTRCov+vzJ3OaoQrdw9SRRJhR4kFA8/Y79OUUAx
n0bGfndTHLzC3m3X4fBWBOuW53oyGaM6lcLTqAi8U9ybDIo9X6LaYfS5dLsI4lar4TncGFAqGnzn
ooL3hR2jzTXCZ7NnJK8iV8KeBR2H7dIkWDX4j1d7CFrFZLVbGN/OjrZq6qn3yK7oSU+QZQJt5QxY
zOQH8IxI2bvImIFQMylHmR07Az/wOtFkV9m6sWHbwtrCwKZOf1l4eWe4vKA6NlFPXT+Z4VkPOdYP
+yIvlVDykXsyaz+IAjCeM7PZQydFDmShyjAjYCVL+YuaT+BWxn/YdG4RJ8wA+07gNJf7ZSglwMG0
7qPNEla9QwSkeQ9hS1KDG7PSXZvGQB2fLwY5otxR5lxY10jU3Aj2Z8otWm3oq6/TWuabOHEZLG7E
cvRJw/pKIeasjRBCGfk5TzHHfiZ/WXcM+dQ2izCsC/epF6TnOreFWiLsdYh/sMSJbwiCdxqmTjbL
WkSB3Bm82VXW1kar5KtquniR70wnwlLq6MeIq1J4+BgGoLk/lLZpdD/QcBtlBd0geKZNTvSDZCOD
ueNgJhs6H40Wq4z0fR52eI4anRrxs11cC7VH+Y5D0L92j7nms35WoyQrA7oxtHMdWvOH4xEoeqJZ
/X2fFcXsa0mGM5wOFpZpLv3OqRvJEA1F+5lMkhtSY8qtXKZbVXiM5DaffVjoz+gfYrktSDIgfCPN
vqWr13CuYcF+9vj0Lby6S8pqoUV58L7GD2CY5D2Ai4ahfEXvn1uD68VmV4ddRLGLb/FR16hyOx9K
vABThkXwUAhsCDNKQI+QZws8WGox1ndaSFz603sBmwLlMfwTgRDPnBvVX1iZ017aBOqxAsySpq41
+MNe1FLM1pucg3fWVmbOA1j/Aw5/5lLLeZklsdVvio+YP3+PeQ2SWeUwWJVTCjAU1InnQ5ejTX7S
3x1LUHxyVHB7ao8d1TxnZ6JRAl8bXn6V/HXHbfC4WCaNOiK4LKQzs+4SyMRuejazMfwehH3gsJaN
F9rhh09wVhq8njE8ltdNLkAqklOR5XAeb5DnTW28uq42dCP6isjycORoh15Oa/dEsAWds6N5sqGi
FeX6/FjlT9JNB729Hna9EXnbkQrRKKBtpW6yr3N6WGS+owPMCt9/tWQM+/QGExabOD8NUrNRRS0U
ETSg3pUygsN5OK18Yds2KMVAVZdJlE4wee3GHsxKDkwyWRzemoDb4lD3DwBgk+mWlwY5CXYqMRnI
nhR1g/X/lT18wzhMzffzshT9IdkIeywzYknsk25whHNVNzVgp6WDAd4WxJhgMaP9ZDrU+eEVrKQU
c9HNG01pG8kP54NOvjUyRkAXoRAvmKw3mpCd6vtb8uvrGkaCzWVwvEg/Tf3piT97ZhYkWIGAGdj8
Ii+DsD/VL9q0aUcElCVl1fLggrSpJLU2OzrCw9e58xXPFYiPyeK8o6CfUPL3Mv+SuHsWQeONHPZy
6rznH5dC7/3IQUJ3DyeQ+4ejoqfHxFFFQBt66VyObHqBmm/rfaxBYcX+7wKBk0C7ivDwWV6QiQSf
vUnPZvjPgsQCNIjyWR/ymNAxUD+5r4PcivXUz6rutF6tlQQ3RpaJuQmm5RtWFhBjQQIVjnmbq2bv
hNP+CW4x80RLy5epfOftThr5nAdXRsIc4ppS2beCkwmSdGjHwuaOzBIIZ+bPPKf6jI7jm7o9OJ9G
WlevgSJrPXP4oQ+S2NL1U33tGhO0xeiuIkzvC1KoIIyE+QThadnMJU7sZR6lQajqrdl87P9G+rZr
PZNYxp2XWxYyya4GtUbD/QPR6fhv3Y8kgct8/7bivoOpQ0D5NPrfBxTGBAXJSUXupvFgzFo97H8b
c3xvgsjiP2nV+REGOQXilbPxcjDvkeHOqCvwxUgLmWyHmIfL5jm/Ho6hssWqf06h63NGtFPz4exa
Lfmxr+5xSv+2E6Og9EAzdTN9mc36zK731eACfeQq6oi4zHVQAOki19TO+dtrP1EIH37vJ09pqUb3
hIw5wCM3oa8nPKtKEMhB0B7CZeyP9rAnxlfRvbaQWwkeWfAX/bAcR/5dB/gfZTcbCEi7SBUz5Cm5
8Abcw4fmRd1fo+u/5LSESJp5OaKkeT8Ta0EQnV4KqzN3fFvl9k63IfXcHnfRrbPU0pE18IMEYpDH
Gs8LPwHJv3t5ToClK842qwp/2H2Sk69BEUHWo6OB5K0mpDojUtUDkZZJGrugey8rKq9rjkHW3ZtB
FuazPzr94T5hyPs014i33GsVlqZqLgMcHCACbbaFvp4vh2JCz//0F/KBXBamdZH0bkHiLH5q205S
WiMfTPjNs7YjR+m+3EMxtCFPQbZuzxpu0ORRY232FHU+SdUoknvT0Gjg5w1B4iupJ7jQYkJFeKWP
Q0o8Lx77o9gFRTMYsQoxs5/QqjXkwOnsE3IMuP1eYW0ZGEU5CThxmH9JUFUYzka9llKvHedxBY3S
uGSsd0p7EfpEN8J5UaOH3aH5QaVHs6muwrO8BcNO1UcgYH/UN45iCO2spyoVAOsAwr+EIn8lvBVw
/SEqW5wdCmf31X68VpT3vbx8txeVRNArlYksg3+OByqKV+EDnIiitXdCOX/m8FJsthFOrgc22S0c
MjOwWE2zv+v70hYQKb8nR2HWOseY4ZEb9b3Mttp5zhpFFKah+RUrNjbg9H9hGijrzTygXhwW+GtR
U7fb89T+GipwsxOYs1ZnpJ8SnkjykN6M9nzkeB/hSK9+6k57owIKniedFjlJFodNbWdPz6MUR1r5
CSzqhMxlDWJ6AakpqgxpuT0jy1SGcskVtuZ1ADN/XeBVA6IAFEljVlc2XjVvpuTPiQs8sMN15+re
yHSnPiJ69HhXo8l7hFwSYNKZz+7SScjYeWetS8Y1NkYVgj+0CrYwH8iL1mU6o7lasW3njBzms22H
z1EH4GTBBow9spcxme/WI9AB6TIZie8oayggGSLb7A5KOfyeA52SL1wrspEj/aojFtHkfhFAIj/H
OVErUp8W1H1BIEdE4fBlFJwfj/Xe7UGr2gveXVDbIndozIC28hvg/xW3ISdqIriIA7gY8lRvK9Cl
EUO0NZqsXY6CI5OEjXxuwujEzdjJPY3UFCSOjyqL7s3W5SkOq9WR0F5w0krcWQeZZCEo2K7hxWOS
dS6N1HUMVza4aSCL1fnKFFWMyP/R6/y5PfSVtqSOAAL9Hx9hP/g+RIyv1AfJJ2YFsl7s4K/Sfcpl
dUFKIBq81qrxUPDUf0xR7ceBm2g4HTbjOtGFgrOqA2EYNz1nRiaDFXAhNC/91k02AIFds7skmnOz
Xs24JIr2ZpJ38nT8itxOE8f/oGfSfTEQW9erhEDqOo6F7CFz4k3q3xbfypAKsMR5g+6gJBTa35Qj
ngG1Ab10YPy+gvm17gLaRcxtAJjp8rmTcWHGMk2pyilotIwz+7fc/yAKpg0Iu2Uo9xDY50juUk3h
wgRVE321dG0+KIqmHEAJhvzY72cFSdGDSqgVpCzY3NhNfHz7LZ/T9WQaSniFakIz37JoMPbncGUg
RWtVadyA9y8cOqiyJ45S5pyS2JF1KZjfqASfYfLyMHl3aqUrpvWF51lSr5KIsVSBbFS/F/QRzmAE
1AvSC9CwUSgzvnyAiCwj2d9YUkLp7sorsnp+oKPL8wzbeVSim2RytiAJR31Z4VyXTahD//+xMK4R
f2OYdD2AYzxpr6uy8HVSTVBlBvTnSFJSTqZIxon2WGbEsnrXO1p5I+RShy7kUtdUiaSxuuL3dOuB
eGthkMmX0Gc4/mcPrnt1rFtoNw6XHRiWNMluzt+D00L83w8KKFl+tLN/hJwzx2vQYJdNV4iwVhYe
O04Gp/jF1Ly3JimtZ9FTfqyYed7Z2PCoGl2zWQHVy7d+rovm9Qo0UJ+iOO3nPDXGSaHv6DNrACxt
IXtmRAbvG38nOXNlCbffqwU4K2v7955tbsLWi72+QQcml0HOUAj/bbp4iQ5tDrF8rZy0I354uJvq
MDr6TmsVMGfjygrBcj4TuLzD9EE3zOvNnBOANbyeo5l0EXZ8KSVuwkAXYQsKrGpd/YgbHnc7ls92
+NGD9TM+wJuz0Ht0+ZAz53zfPwezPrP4UDCH9jUZ7PqoNaCQkQJ2Uc9gS7s52Pk7GVIFJm4qFUMI
tCwaNUiLmRzLQiDaHz7/wV8JxwQkZUMQH/Or5fn6dga3rgVVwdMD8nCbmcA0+u03Z/z5XXVccIp0
/pkFYVgLPSavQwxRidrl2zsLPt2dxngReqX+12Rk7na/4DEe6vPrG0YJ54JsANlgSDzYrhMbu2t2
a0H9KAtDxAOaibG2AH07mGHNJ83bpvGTS8Yx/y9S5F8Oh2UFkhebHqjR5koOOm2lxNtCOGd/vxvd
x7+wgDZnxO0QJaO5XsiinZVtjZMWnCHgPxlxoED/gNG8UXe8wvPtDgL0tT+bcZ+rzL4FHNrhEiwV
hgOXFocIt4jrGmNTcqcYmeLy+kNcPfdZTm2Lpr6eL3OH59reh2N+l9Ytvd/jRQcs5IAsRa+efkgj
MvrpWxUuVufIuQrIPXHrr+j5zVK/D4gyIagRNnKpK2HfWlBWqrI+wQMu8ZyXENQMjoZH8g03+BL0
sncUqjvHi0Wz3hd/ZEAtfi7HxjLL6Hec1pkEsV4bm8ZTf5W9jvN+7cxTCVv8ZYoiji2VP+6YY2V7
zYv7HqLoNt2IM2ES4BCWFKxTfVg245WXzRY+cwbTTMNC5KZ5wSJLVZzVMSs6SP9MEFVsOLoAbtIV
PATGehHr3qMIUcU8TBTBQ0WTa03b5gtQFKDNy6PsiCe+XrvzpTBFiAJ04jh1J/kOKl9cMZqmiCjx
eVaazXEImbQVBusJNQiFAvIUByw6KZnLogqKHJ4tz3YxIJb2Woaukk7rTx8qLQIiISzJ4JtTrJMi
ivxLTvoMBxsUwTHU1YaCW2FfruaBue/fG7bA5g09482nDjJLUzftFM691VS7MSBKYZvhSEsgiGZp
Csa8bpwuP/VD8lU5GD5YPWWkGfaUtxNVZTOLRMaExR1cnu0JZEnH4gOFGuNNMveN9hj6q1AX9kUx
ifqbnk8RKfUkVvvLseMC0uQhZlIjjVDfwIxBgD0n6RKN2dlGxbGPu4Rc9ete83MQU0zMRXGchEvg
vcTT2jpP2+pPdsUOIpFTvb6yeCERISApDU7/Uf1yfnBAEKoYOFu3RfHmM1A1yByYiyH/ueTQ16nr
cOvKGQAja2pAGKZov/l9CYSksccJkOrgTMx40icu1bK9fAHMJMNvrMN1qw7RegBrCa342lIupaZ9
rqt9Of9wxnY5SjsP3vRjidtq5XYIpWEYFjaArtX5a1Sia8G/+C9n/ZPxlkKn2zjQ0/+UJaLQTaHy
PQztecTVaXWugjWYtcyRA622SdAEg6/FrlRft5cd6oA9OC+SFE52GlUadnnFR5paGHGhAkuFE7zu
dFcEUi+oXrKXzl02yT0Gw+zV974NIphEgGGRjL2B7RnmJkTkhUHRW+TstDRSq5v5fyzLJXZCBbC1
bOvIsDaw6Go9fAySOrKz9KwVaRLHJMp0G5OnB60RIWCPkxv5RxBttrJFZROcTTrCjlvrYoTPn0lR
ZXKQWZDyfs7OxGoEFGHsLBS6DQLR+8I5H3F6bEHu/jTuZV2/QO63GT5/cVYSlNNtVE7SudyWIQwN
sA7mf54CJ/kMT3O3UCSXl7mmsEFKcJRpNc+Dlqj68SGWFYzkZ+PDCSSw24yXNbGEqoyI5JUeV3tM
wWUww1PZnoNjINjtXqM19+Ci5SJfQKEs2sE2g4xzROAEx81NY8cP72TnsUTwiQ2n6s1uELNJiVJZ
A6akW5FvLPU8QhCX6OJx43sb0LgZnamMFDzYL83Y69+sAs1mt2VkR+lkM056DsTN9CJFJxmjanBu
+I9CxSu/K7uuPd3qXfvFzP5ITqdWwIDBxnvcPaQlLIyKzrXDOCnyzMiJSogTP9hHzmqG1/kOS1o2
hATXFw7oYIQ78//XJkJG8qCuiz1macLBJj1mpCmH3whPzQPKjnlHs+E7+4NO9WgUsFG8wER6AJcN
c8tg8cI9IVbAAcVrV+e4Z3cOUVbJT3cA0z6FC4gUn4RUda0UV4mXb+9BqQ187vjTVYKK5XfJz/YF
+vX7nnTbvQIsO1v/i3sDAfK4VIQrZPZL9e9KoymgNMOxGXWWMGKvIuxrNfB2KcoWqS+CCBPDqQ86
mju0llHteU7HH87IocCkw+LFXqTHKj0dxR5rDM5cK5hvqMspB0EE5Y+5NBlykQky5UcisOJcuqGi
bosYVUnLjPzv7f825eFYtjs6mlahPQvVigmLQB561SJTl5+G1Qzk9vzEVumB4X2miGRxDrWpSxRe
91tYtehG5BKAleHivXs6LaWSyvtH5gJTOYQHl7TD3JneyduATBj2a9TpuMQvGvhLeNrdABYlEF9i
EoqjlEUsyfa2prAJIeBcTcg0I16miJCTLDFSjt2+h4bcCOnrJ99/HWP0VPQEinJ6jSVg5loRd+so
Q8VjQljFnbuJV60EKAIkRAk9QQNeFM3MIq1ko1/5+D8wZK34rbw31eaCyO1wZLocBBoL6AbgTaIT
HMfamkF6Wh9pesOHrJlUtVcNvCLHV2kJWiSaf2zXQSsTiftdEvWKqhGrSLSQLi+s8fMFX6P+ms/l
Al7ozK/BAauyict8B5jq0XIIWxQiWMbvp77M/yY2wL/9V3WfMW6FhBYqP5xKr0FsrpPw0JokTf6O
tmrPudgAsueEVDDLgKXSPfBdVFrYat3tLWzT5PkT/4eqx3+YGvYDHNYD3JMsrmrRjiXe7qVps6rk
RKvPxMR176kXPxpOopDHTteyQKUVQ0HiFP7TGukdlI+FXFl7H4N9LCTzEBviYndfQ45nsEtPs/ST
o9gMQDMKAyU5AUaMoXphftc9aowZZwZw5SyFZmT0V4micfg6esI0pcZ0SUbwZcPgSNCgxJ9Q71D9
1Mj2kVgxX5+Vp4KK6JIuOgd+QoBEddDU6acVZr+stTGOgkZn5bNsMaXpnSmVfxm9wV2YA3QH5/Tq
SNIg7oWwYy/++Vwg+i9XkCmDjfnHqSXtjcViy+HkbJlBIjVHg3iOjGTIfpgajFKId2UzRV7ygIhs
vriCC9P4igJbaJGZdfn1e+W+9T424puwyUenwYhAQ0ke2xJEdR6ejEFbKpGSfskQBR5S6I3GzZQf
gW2IIyMhgEypBzwEWaRuCE5PADKpB6bHGjqcC/xuxFd5SsM7DI5C6lvagaDIUpi4zhXTa4knxoQf
CTBdd6trIlkp8zGvee0MKZY44knKPyVIbPFiN8veb+02S+xzdGxnNEDUHDgMetSQ7eC4aBe/IQth
6dGjz6LppUqfP0k3DkfmYppdj3+mYg14LH2QPYsWi7e9+7g6fmMkybymT7O3jmi1DdRq1FSGGMYA
6dmIOKVyGSOrQsNU3Ov0kUYM7lg1gyO9+4jg50EeAd7gFwESods8yfpUWD9IIU2V2kJStA8UUEQd
84imFk7KUNvVKQXimnDdD8BWRjrFyyBYTsqU6p6i/JHBr3FkmG8ewZplTHVcmpmDY83BVn9+pWBB
p9+DpJ2QnA6Bn/poUuzjtom3R9rmLS5Nm6W4j6I1pNerIGI328jubdSlS/IyfiJs8AZeU4Hx4hq0
EPI8yJ64/WjpPqiSQSjelVL5+SUBgT6DG3AugeHV416SAwtMGfcBLT8EZzUltNlXmYTtufDHMguT
cZ+1WOhy2m4yaZCaMzbG5Ml9Bm03YEz+EaBAbFYBkDDquBKW563B7S+EL7M4WRnr/Dbc4piHn4rq
0ULSbFcm7LXky7FYtljCYaLtgfM6tjcGG5sTlL+q7qedczLAOf0Sz/XfWuf6we3k27vRmEdOByhg
GbJxBsQcGUSQFB/nsg6iCRl8vA0j2I6RykMuMt0ZVJAFagrQi+nOdXgK3r3xGpk4hzv6cRZp06DU
FxjXL2Q9aA5TAH6T84SUWAbAJEt87J/xBWZGWlqHTnZb5xqwQ+rN8Qp2klG7O28RBOw6JzO7G+kU
7nP0tytIItdn2MTee1Oxg7B8EXUoALamgPkzhtXNnvic3raImWgfHVRDaSpIUHyDxYKbzqT5Rs0E
DAe0ZNbbma/8zhhSQMtCEHzsOXA/LkVIQr8ZPgwMvY6R7WnRSzjAiVnz5Y28TemVo2Xt/5rjlWXs
T+B7EznMiKMy3i+RG2tzsodPwFE6dh5mkhpFIVLX6C0886Zfh8Hm9nUDN4zJbgi4vSzRLeixBhoQ
WACKzxDftcMgyXR1bSV02a3DZv46f2WI+vYMspx0dCOuVCPNeJh5L0BTh38uLBrbkTNB1qbpOSfc
ewAZdR5LbjBY7LvGOkPGj4Hq7Ki4sOW0Z0S7YI/MjhS28fgUqFVMIz40FQop5rnIMP/TrakL+Td5
ZPlLaCaVmCeqKW4cnd9OpKh1nw0bqoRY3xtz/dy8xU3mFmg5hxMF0xTA9XlkvtXqamtK2uwylKNb
TbLGAdaIT4Ms6Pysv29VRCwFHOv5Vw6WYuof/6NgYAh7Z6/MTE/n4h1h8cHwvcGgNYUcJeLoVHN9
XyWWMcMZ2QvoQUkbxtEu1JyYNyKpsitZUVzE1E2oT5gvdR3tdyIu53tgiQ/kw7+R0BGK/Vz5crBl
cw3Y/YIQAjEgR1y+M/Ebs0YzaOUJ50orn/dpcG+l04LKdoE43PvJ8gcLzNMSPMV40MS6i+Cd6yD2
IggXqhUJt8FrWysa5EaptGgaV5aArMD7Q2Vne+nZ4mVo2Rg0zbzhXoXcOdJOyMqYhAVNb7kuWPdl
GthgogDzn0BhBi5h5M3fHucCpqNSff2S9Q44engL22gvDpIKzxnSD6Rwd8c3owolyVIMIwkKvncH
IKX4Zg+aEs/1UejbL3j71vhmfWwptJExwjjg95Hh0WZehjMCoCVuw3Z2jgDGzwM7b5biqbxD/auC
Bb8knFkP48jsNPz7xlHU6lj8+xhVoU/roKT7fr4mS2bS1cGUmD6tBiNummBGLGz511iybTvr79yK
94c/tB2QEBAqtUdG6aJ8GXpIZEXVa1GOnZ3/mTYK5ReY5v33+X5fHaBNf6pg0h3rp4OQ0LUvD0pb
Yt59N5lUV6L5DUDKcVCYwhgJy8mQb/e9mNKv97amLqfImCcYhqzdZNYJ8rZSiCApBwe2UVsuSUqb
O627zQQ4v3GpDb3DYnBFMhUJZi/f5Tcn9Ok2cav+PIjdqpI3Ew4dSzSqbt6qvFbr909o8PaeYaux
5noZjKnuoB/ftP12vDt68EpxKV8cBLM9qygpmzjpUb7u4ajtlFoEstkmZwn0S1XLfeHr+Q3kcbhs
OYQAWYz6QKYiCL0uD3YmjwQL9BL3+v+h8d5u/yCiUwSodKR/JaOf0aaTpzi72qZQmHZr4vjb/Wva
/ADTHg/6K3YyQHTeJhkwpid6ME13MsgwoZW0BXmMw1Y6ll6RqfELT7SVP6h9e5lvLdOokeUn3cYB
+WamrLlPXc4zMwjuaMKdPSU9sFonmxTFqguQpjrQwcu9aJYVboLBm6JA5zmi3wbtoqx1tz7Xu7ze
NIM0buP+zfjVRBu8YSGKmhN5I6LpCnrsb1XuaqT57WP8TARBLdYMvLLfMfrvCl+/i+sMPjA3WLlv
vmwt6NYzOhKAbvE+y34QaEY4MorsGITCZM1k0+VwrrmfPFCn5WJ5hC4UXqNXC/FpMzFkw1zZ77YO
hXTyLsLmzzFn6L77eKdKHa2G01vsR8sM37DZiH7FB2HtroLSPpeGUqp4M+aKHTvc2x9CACD+Ma4C
Cw1Q2H7eR1pkfcJxyEC0ToLU63mL8Ujyaj+3UyUFAe5WUVAP2apGhrnIP1Xo1CLF+wUitE5OYyl/
nm6v9FJj92zrqxE7MsK7Dn10ktR85S653IQNPfW6BIzV+pTIezS+r4uG8nhJrZ7pPwWrofoWK4fO
BuznwYKVgsN7Lvve/TvnUXC8jSYwOuL+pRnnCDWOerVPKocSRuj4ir8So0gH9+5eDeSKH++6hDWW
5ZfGtKUXcvk/LEQCIA3WZlJq1iaEtp7cxjoLgjf8sb9OAdEwWzwl0nDIxm3MCcWI9c8uxEFYe2I+
npV4tOHSvHvT8mgMO5o1G2nJs0FkKHwF7CeMJ7gsSHaafowpVnU8vOmztwfq8YfGy1X8yOamVQql
S0yq3l3OgU2G58tCzbNeWx6o7zkSK2AP1gMEaBqQlnabyPD56HLRqYQBXiAkC8CHyi4PdM6P0gou
C/ySPqvGEsJNZNJxmjliHI0M+9iHIqSkBaU6/zqdoT1GjKqIwc4d2UP28kZtPpzU75BjP5lHooYX
ZxdT50N6cXOtnHxTC+k5sqBugL6OYWyLRoAgVlSjmNbZfNVTs6PBx5uZfaHCFpx4sBSHMXDHYvw2
aSIAd/+zw6FBnsQ1zP9viNoliKOIUj7rtTAIJ1KEvMIAMx/hkrCwZ09AZCajGAOIJ4FLvDT9Fe3Z
wA9qXaxbIcSjGAlimy0oxYCxo98XMWwWE1oU9PtUgR1F2UCTwS9hYs6Xzz679+ioQIYGJGU9XWa7
WuOQCkmkr2IpjoMzup59Sun+ZaxxK0ONHMyA4beKHr+qXZRHZlaleRQP2psYxUKetgO1ZegQoV1w
uDzP8+ZpYJB0VyLSS7Yt+hiy6RWlUYJSIiInRRGiuwq67F6lp2h2C+75m9+1g2Hrl/Rqo4+ZufQc
Nnebnl+CfCnBmWpeWgSQTl8KeXZNyx/3dtCtOxRe+XE0ivW75ln7vq3gIqiEjj2EWSD+1wZvzSS+
IDcE059M4VpSov/oXtPAbDND/gpbKfo0GcnKS54EnEfVGi+9/AxO8vwV+RBNiRklIwkteaNXAPcz
Hf9jY8x8asq15l4cGpc3hBKpfLQivpvyB2wQLReqihJmHNubhmrSHiOsXxWnv7YsqMFlM3IPQe01
JsUY1rTzjqSNAfKDvyB8qWJxgi8LaQZQT9zDGmWbbjTzdtDfibk9rgiKOdQ70cNOEnMV8O+mH8mP
9k701kQUi+V8wBz9SPsm+lVUJDQrrlvpyYLrRUcYzSSexfC3kGbWtQUf/i1f/8CrZgVOZjvrdclU
hz6f7ofN8ks4Ciew6IHyBzyq4yRmETve8/u/g8PlZ3K7RZ/TkxRn8TtEW5UmdNfwN+/y2ePQODgz
pe/t4m9cqUeluhNiF+B8p4L+rZBIoq5Y/6EB+9PEpf/oxYf7OlPtgPWNngABvP9Uc/0Br41F+Pjs
IsecjmnqjJQeBxDTGhY0kKCnn503DjbU3YGQoLfXtGbkUPlBgi7q9/ZxMY3iJ9nLZQI7oyfROpiz
5RcsP/FW06uVev0PKyjvZtFcnm7LVwhrFM63SvN84aUJdwKWuKqCVgrO4iJIGRlGesI8PScEnW5A
4hjQ+Mhyqk3TXKJJb3Tq6F1JRh1IjpA5xZ2kDNusnU6g8N9QmnQb2MbvdeOcyhH9GXIumIcE/h83
mFidzhm8LO0PENh/pBPE3+JDD/C5ullloqHxaqI3EJgmbx6KYOMwVX2xgahT6jiumFoHJsYysu2q
Ae/+kMeLtWhpGOykvlPgkbyaslwM+l0VO3oIvj5i5mqFS+mSfNDibM/4RS/DDof2pYdVJVJUSBpd
NuRHVh0s52oGQl3+evtsmRmJRP0ShBza8gtxWQEBo+HJb9hsxxV1mAKMnC5X3Vn2qdtyIdAnzxbi
cJt+r4rXfERO0s4D6UVcstnDaxG9tjlr5oA/u0x1NWTGhuKyGmrYfEsMfp4xFlFZvoGoYBR8yBEO
Y3cQGy1Ik5FIQbfAHQoxvT8GCKAOZTAA4tWUems0mtOXbNCj1lttVs3zQFMhYP6eWHtxqGPA+EGx
qrXkT1VJWY+DetCB5dxlG3WlG58GNeNXQ40uu9KKkjJ0DGkimDJO5N33bS7OQVJcWl8gULueXTlV
yXEuazgq0kK3VN6fbEGB7sIKnuRIMyK/e0G7H/Afj0o94EPVniCxy1jS5Pc7AWsb9l2pVJC7ax/o
M4JULY3mUyL/OeCN5AvN6n62nQBFVJU/UJ9WeyjuP2jjMIUB/Hv31FVyDpl9n0FJjgXeR7h0AZL7
7Gr1010SCJAKIZLbAb4+bEHps7Ia4tCzohpOMFXg6Em2XlI3b4ZfCGserTztq3Jv1FFEYQC5fb0+
Echzk23NXzY/eqGktQYoz0bF+33k+L2hE13KETu0nrTkH5UdAMJbeiokIsW+SVB30SHKr+R+Xrcv
okPN7qDqvBbFt8YFKjvJ5cwsfiAkEQsI3799okoAFCOkBTTIpqs3GJMYjEODcsh3wX0sWDMNalek
AZ+jzzaSTh0iNM+9mfq0Nm1Psi5yQOPSRLesE1m8sKlgFe2Uf4UwC7EU8g0rk/UwsYNGuABMny0o
BMMrcQOc7wDYxDLbYYphASYdThVCKE78Q0yKcldLYwzcDo7kmhAH1wLRzd6O7vwIwQ9zi00iGvtT
FiPMPHlkKPod8/CKZoSzMOr/RLKwvJLt6JRkbrsXrzutSsStpLZga7IxsIablUnnuuLQn7cWz5zj
RjWrbs226cmtsegcFkQZyDHNjvS5TQzVfXOByFIOK4jjitf2gYTOTnNlu68SUbt0Z+FIJ2+cOGvB
j46uIty+xVolSthYuddeXk0yY3766AjJoOSouSDptBSKtiFw31CHIEMDeOk/I870LaF0e9XCFFaP
GJSnq5EWbPA0JE7mzOi2DAIHBvhUpOTbsfwG2DPD/JLgWUTPtnwrhbquvOGjhryKdGCIzMw68z1J
w32GTZjwBqngsfDHQMe4sC8WTmthk6hB7NPfWnYZMCKXCdiCP+6O/+usG3CQgQSqXTLrjJ4J9ZbC
HMs7EEQ6kEqRkoTIoDGMRsl52A3/jmUW8SoS7kCWH9xve/IC1txlPRJe1C16MsVWsLl59+3dZLbY
UuBBf4u68A3VC4VTcdIUItI0V1cDmkq9svuvAySe3EoeN/03ehG12OJ82ksj0IjJIDrzmrpbj1VJ
RH6wJvQ3Y442gk98mn6Ir+rAI0l3XQRRwdMYzh+K/e3/AsprRq3o7Q7ovxKySlwzp48YTGNTgADx
srmJA7OzvH8Y6LpXW/omAcrvDnyxi4MaVO3rdAEtoYAX1mhSkiiYc4DgA/mNGp2dY49Id8I+b41y
iLc0dYxV1Y9tCNxmUHupTUWF/lUi9WlgSLdJGuC0X9Wxq2UhjuOxy+wYVx4wvr41dvgKEAcwMVFm
3QMPOE9ni0byGlofqNKaAkPkeJVMeHMlbJMUPuaU1balHu/m7OKjzWHtgdU3pqvgU2j0TUjtGUmC
e69C+ZS5ldiDdNEyqHtscKwK+ry4fARqeSOTO4LDnzXwUcv6Q1wZ80ZK2Dl7/cPgMqdvTRGznd50
TII2EclTuDJGsrrkWnPutlyv1H84x5ck9NBsYbTp/rEKGrmkywfd0i0oWjG4fFecHCCXomgsPqzQ
yzOGzpJF1+4ugt5By+DhQSMR1dflMN4bI83/T/uTy5h52dWpJopvmzHhe6htFC7C6/C9iElJ3h/a
WPPpd0F6+j6Rd8SxdY4adiul4FJGtwjk16A8Hk6WIGN8d5phXqNK2pgvsut1v/z2bkZtU2tohq5q
ONDnYxag4GegKIZZjWcPYe4BYdGRqhlphFv24B90NecRcbB0GBLW2S3b+NPsjjQPhBBrmRJx9aWM
OS0Wcda/g7W9PlGd6jbh2VTsTbqDhe/j+GPXF+0GtRKvjH8WZG11Rsx9oMo9ADMhYQPPgozkOBvl
VDMSBuXijDAj+dJg4HIu4JtMiOg4HJaf9uzeDE7q7OSWaN8rFBT/5lkJS62ME9JvjEutMxo0rbkV
te1eSDcHRu8A98/momHcesHjHgIX4u3+yaH4n2BydFsA1vft1Xa/71q9XN9/KBO//StBjaUwqU9n
TjPjnw75cJjcimi52naE6XYHxIqxFGxgpvvGNQc4wDQ3JeEFjqY1gq5RZQieaiVlnTivURR1G5EI
2ZRtd7huGZNmuR0ySsOADWGHg5cI2REMwfyDEsC62PYkzTunQGf2h/PO9R/ReJGAox3kaaO6R/EZ
bOvhpO9l0LPXCiXeyDt/FFuV02lIO3k56n00Ksxj9MNKWMb5jy+IhP3Hcgjcj+zhKGrmBtbL1ed4
hagbsa/AgTqzG4YfOg03q0/yqLRpouE7XcvVMtmhScTJsZLZKLgBnLX3iw/s5DxmbawYY1e3YpMU
8vPufoQpGJDQ+gxwRKUlg2C0AFKAULZglAZGYnS1wZ79gjEgrBNZWuFtk27PxDfe6c/Nk4eyrhaU
40Buzg813TNAjlegczopRlKKXU8dQQUEyJgUKXQh6y0TEsKIpK7VLynfB4aRn8OFvFJbMqEguHxY
MzW7zcD4vltnqwkv9r2mYg3ihPgMB8LvThtdmTp5gq2sxrzwDmcaIUf6/pq0EDizSB5J6+9v56QI
2g8rTWaWVGgg8M/x/Ktw4+jiJ+vBDlfVDFM5/sFEMJI2DTkN5QEUFHGNljx2Hon6E3b9TfR2RgnJ
lHmBLafmVly89m3vCFnIW9Yt9v+xTfoXRNmDzaf3Yg1ruGFTvaNX2p1SFBrXGAvtajgKcboOkcPh
/RFwFB/qdnTPGzX9H6njAg8N2/wfDetWqMNzuEtUliie6xA3g9hzSVDvkr66DE2P71H51Y5zapiD
7aG08rrooaRZYRnAqYbWXZQXIAXNFrQ4FfGbDSlG4777dDJVahDYGNZH26/z9fMGo/Ue+GZRTIAm
zJZiFJyFBQPt0P1NGBXHljxClAp7CQsqNpjeT9IYcoBfNjavdcV34sn+IN8MgdKfxFgKhlbbntwl
oa7gEfSnSSNKk8egIhFSgeGV6UIh09F/y6DitDsXXijZBy9ii7HoiLDjnLS94uoweHm2jPZMfsOK
FipfFqt712JmkCgjjU6/V95wvXbQF27m0Tu+0BLkviuOqB2mFUUWeBVAzY6IGkImR5UuPE88RIks
YOps/1saP5scK2LFvxlROvBg+7cO36h1bYbguc1Xjlp/3hFOa8ddVy2z2rD0QqF1Syz4YIHURe0O
ZRcd8HZGpSo7a3+B+ubNnrCQxP5oLHdhSXFmrcq369jYqGWAnLQTZUyg9V0KakWsKfIaD04O8zeK
o3jcrJBu1N3zcqv+IRUOUotrtoiHk2CLSFXgLJ9IU1Ajbw75A8kJSqBUH7dgfCVWAxYqeBnZSO4r
KVG7soAMFrs9txQh7wAwvg4ibRJZDoldELt/c0JDRQU1lpAppYDbKBVX7UO6EGF9NdMwnkiB/7/R
5/8M6cQf6t01t4a2hmfNO3P/sbWOkj2JDbXuxBfJTQxExfli6djUO0bC0vHNKHBl9jKeaJZD00Ht
vkhTLe/g0AwKyhQjYD5fazvPCxMaVPiAqG2zs7a/2zti+8tO0t04w8fbRUwN4+f58Q99zHQvwt0c
T/46WoDNUXzEYt4LQ+Uyt9VCa0lVTuaBk/ulYTc1ZUIoVy3yl1stPuMUMSKWV+U0XQeHFUdpTvbE
lDZEYyV3SzxI9N4JJJ9raNiMXbUJfPtdgmvjKhYT4Wqe7+dUEHyYnoFqALeXLPsVw5xouekKVSOH
/H7pU1BkjsKRP/pKMHWlN+NQiXJs2btqcEEWujntrY8wqN8DD/JH45+41SNqf/kB73lPHDyUPS/T
SVxqU4yeES6proJdztb4WLxuTdmpQ1GlFfv3GEsuEmI9alxc1o6ku1un0gUvWFbL0g2Zjbl2LLsa
Ki+q/hRO1gR2zLp19zRoKVbyrVMiZvl+zLiLoLxhDPaStaK94YLaX9HHex2qjZjvx8JKQMFfx/66
sx7H1wlrqHM0eONZE1136MIOtpiDukaLqscWPtLRyMA8HJuNlluhOBoX807gkxX6XqfroguOOspe
NbWcsvmHyAeRP8cH2VPxW3INiMYT8lbQmspeDRntoWD1g/+JvdaGHmpTqpX3eFND5RL3y+/i3obL
q3EDd3CEGxw5dshGXpjf8N7WcryZKQzYvEETwTdMAW1QIpXcPeOhy1bJfPUOuWO1tY574Vbr1WXm
vngQxg4A7supCbSBbuhSWeO3mhgKa1ydmo6wLe50TqBa3NwJvPAuPQ7X+T6aiJ69MwMyo4rRLj6Q
JCFVHHXflqxnttMPnIBLRKy+/O9C66vyBpM1i4voOzCtiC2tsqsMy7wklMkkYlzsrRIysZNHFD7v
Nm0pbZPM2qJ340pt83wTp+kMVX6fSmt7CLuzVc2FwX4AEMJWd6g3Z8jev6ttiE1qQbd8anBSyjLy
flfXHVqcrcCPVrqLOnDfMKb6OCJ1aaiEDrT6hCz/XKCKfQemEyQL9QbVJ2RBI1SCeGdnwDtslsM1
sq1xESgmVVac8sJaWzC4JCdqrUx3qpAtuoV58BJdF9pA9A8fouOwdY3zDJQ90A7ParWYximy7KQG
vDm4hLrlVzmuzUh7bOiQTHhzaLfXMOzNm4p1opvi7r91m6yV7EWVZf1MHYDMA21fnRBEA+gwfJwE
GS4zUS2p8Cix3wprkEQ4KbsPB8Tl4JhD1ndGJwCT1Bue84PuMLEmNVZDxTYWCjJNZ/Lr8o2wkyZt
2IERRLD3DmWyvODdiBhi8Dxl9v1B0N61MwgzDanbnW1SM4tJ2wiD6gBYOmTBKuZoOdp9rrBD94u2
caFNR0tH7COfrVMZxsNVVL/69ay1gG9EZ/8tBfiCNg0KlSe/CbAokBMHFi16ceiO0YOed6vDzVEv
KY6iosKR9OomMRFSOnSOz0ZTzD18RlBCDjRgm95QZiPs90Pkl568a4G1bXOY3Zhyx+c+5Ru+fnLd
IxYn98OtdY5mw46RwKVFZbHn0Jd9xAux79b0qCVFmHMOGZVKOzPFEQBJM6j+ufKkv7ikLZ3+03Ck
+v8osoPcS4vHs3a/LpBHbCTikmCWpnllyWPjXZCuvnISTZkYLmayI+jlzlvRHHrhr+WleS5z6O0y
iH7IduOCLa4KY0GtD5jBjOUfhFZ/ezN8O/bS4Zx8pw8rtCy1rycURL4BmiSVoPl1poMfPfd4SdjF
eqZfzVsSnn2Z0nyvtj5/godq5Rbrnjjro7QQrGLnSwsfuM8tPBAmjUxeOc/Iokw4+JWyTra68WlV
mVqzHApdnaXKXcpKrvaZVFI9olhkDobk8wZYt59k+8j/QPBT5qxsky4aJmQgvFRPOBfxbuDjK1h4
c5DBJ8hnzkBuDXrPD3lQgVKaotVOkAK8laZ2kSwQQmDnptFfDFx4AJqQ0jSte650NcZqRCGr/ob/
JOaRBIsV2rzffjU0ky2xWphPEGPLxGIyyCd8mznxDspauQW7oY2SFcb0S7jND1aBZ9IJ+JGlnjW6
fgm7ylLoatiWuU3JVCTvc9/VvLUxKHbJxzTf16Zuuqk1jD9OWPVCs4nOTKdaSgWp4wbeBfAHuFhj
2pLt4o1iqGgLlazfu3vcCSBUOFn7kpBtopqmmgH6n/iiiU6sKzh52TwIcXAIqm3i20jPKuhXKp0f
0hgI8uw+sy6QSoOLn/60/4Jftdm53TyamuhSwbOdVxSGKmaI561+PNi4N+iIhK+aLBIZgM+Y0QTW
NTDr6qMCYKB+hzqA+gWrjoXZS0V+i3QVNvOv3+ctzBPF1aKp8F+gqkIUkHobyMZvuNtZNLrbJGIl
4DDV4TOSiU4eP94L0P9rGZ0cMaCh6wMJdct6d9FQTbHzH8As1AU7xD3tJQAdpzYXASPVsR4gUjP3
kfSYoFTDh18XOWIGpzqOqsHgsgmX3ZrusXZohS9ed+tDJF2AY06qHeG30Y2keWjTp4JDpXsDwLqR
WAl5Lncuogpki01sfM7ffK10deUrxWpMkgs91Gp2t77OnLJmgWXYbwHDeeo0iGaLuvtE6/J71f5q
YcjDgkfOb9q3r1iT61BxSa4iV3f1x4muGohwNcpX3ub4hVc4N+LCN27/alk2pRj6SwSUMw4w+JSr
P71e/t0VCmtZeUXhtvKnIXsfSK/0wBuNL9R4IxwnIX74WZ9OPCJhzMNMCGTye99lCnIBHon8xLK8
Zt+W5+4RJBgq9qUcInmwlo64nbqGVqHMpjsfgtcYd3j5W7eOs35GQ5nVr1a+v4cUthCla9Ld4enS
na1qJ2ydVT0TndkK6rq3EjUvtP/njhXL85AgPrXEoaSuPj7qmyE4KgN8JM/Tsr3jIBbC0DMxbMkL
KYJBo/mCXM2AnckLQtu7lrLvB6KWlydues7hieJRZc3iF65I2mMSezHV0NkSNRQD+zWanyK0l0Nm
Hpfz/3vWKc0lDJnwcG+Knh+nRm3QzT4RGjRV8M0PrCKpK40jPhquo2fMf5N/jTVWwzDKJ5yg72yR
S6hiVF+sZQZenwJP/7mVXMDt7UGk7PLeYdgZwTojXJeYA8B/dan36a8OSDOV5QtygFBspp5DBDE5
byyHuZ9IPZT/CreYQKxvehK5E7BShcwfia2GtlbSk2UoUhEvma78yFzASAoVAUN0KS+m87Bv4pJt
bvPv0NVCdv/nNI374pNNejmDgkwVOp75lUhPKbp6NdQJ02+NAXlTIPc05rfX2KniTUIZLoGISSrn
Gwww69vPN0MBoCi1DpVSVP8h9M8UDdKbc1bBcdcKE4Bm0KwQDgRFp6GHA/Z9ANY1/VaMsDXTdbEp
utx9A3sQ9EJu8hsG2Z4JJFagH6gOacMxOtrdV9sj+M2EjhWgn1NKcWqmm5dkgLmVY+PlAP8Ogruh
sCV2KaBJ1j7jznbn3Kd1TEldrBd+pEuem3JoDFiVqKRb3qP3dKy4jKY3rafMLWidKUpco8q7uqUU
FTqS6BfFaeISV1gflfM4cI2OBOX5hpdYA2KYms39o+GPKpIs9tEuaF/ynVqSquvIlugr77yzm9vu
O4v4+fLYtR4Z19bymdl6I+Gljh7PmJ1CZGD2xNyh723qs2FZV0ne0u16biskyTrZIhpei9UDtlMP
fdW8TD6cC72UqehUIbW7phyd3gK2oD5xpk3fzfK5APlP3PYoVnfKqRrAFOTuSXkaFX1SLce9MKP6
0kk2JMPgabAXcqEEo1V6I45J93ldfJoCFYtZLwwCeVg8SiIUJUz9qM71m1jFQCQXT/Q+lcriDARh
MARFI+t1b7wY0LSPjOFQ4eSnGjP6r5bRr3Q0udvE4ljiL9TOPRHLKW6Atw82xjsChzvw8OVXOl5O
FPXcUSJHbi4W01QftnWrkbcCMJKvIW7Xv0TNG0XTBYUysylxV6f8pyVnE+C6BICy0zFRcv6irWk3
ts1B6LpQJeHMMtGRj0b8XgE+0rE7003ec/knvwOabFCacxguvglKqf94hEvJJfynQtl2cycg0Qau
2Oq8lm2DsY/k2iCfQ1DmsD1YCSts8/nBkyd/kIzYZHEA8XONc2q6y/OplPFDbID/ARZCjHBNyQ0F
vqddZUkM/9ds/JiDPTFNO041MZvjxTDYWDuE42ICmyc/JycviBRMBKY1WMRWI7kNrgMVTI1mGvXg
fX4/q2j/7ck2b34Of0OfprZ8PsVY5Yg8VOWZTFPgpOgb7cTkRItVxuEs/UmO8bzy/DKrBypyEz6S
JT5bGxYPHf6vAD+OpZ4gP6shcgYT6KtxvtrQo0IOGHGZfIC4dLIa0zSEZdVAKITTkTAfsajKgklI
j8+MOdplLN07fBHFr/GYOeDSrFr7gBnhshkIBK7EZvqtwV5uEt2eCjwZlntKbmFwTEW3MRVQTxmP
1fQQmtMro4pTxTJF/aBrZqCXe2ENg6tcoSV94IQM48nu3Z8Lm3+sv2vIdobluxE2r09PP7Cl2C+y
x0Ji+uTCfUfJTpX5Q10tg8Oiz7TV5gjEKPKLovfRtHbsA0JPa6Soat7JwXQFca5SB/nlScfe976c
XLXeCDg6A6KQVLETlTc0TwiOiu0y36g4aRHmhOszsnMydvlLtH3C5Ifa34x1wyT2Pxkq++MRDQ4g
+Ap9GW3wQLcDsGkLYAUXt4XhUzaeS5zhUFiQ8F2GiEcrKxFIIoLqODRri7U1p5pNNgLQkmTqQBFs
8WVtwNpygH2auFXxMv8iPbPFzgDq5tiPcxGJH9WaPTJ7cBAqyFoF1UMKh8+OtRWaRAtpEG2HnV6A
9fBGecccBLIu7BMSPoepZnMAVZa/L2Fkfs+DYno/scolcvcSmVjtlUGtM0C06KP3DA2SxE49sAwe
NlSbgOJUa2wRvecnlYgdcG/6ZCRKl3Lf01/FbL9q7PjkAFWYOo16jaD6ed6UgCODL1ED0/yH6o2D
c5GhFmKZ2wXn2WCN1msy+CTL894XJ0Zhq09Dw9IU7izymgusOThWKv9wjf2Rf6hDZs1Wy0OoSyfA
joSwtyclz9XY/hirRy+PDAGubZIHSnxcK/4xTqNNFLe6qLdipLZgxwmxRZRo3TAorwjj5Xvl4kKT
JbcrM+RUkBHOCiWvf6r/CZH84nL12tRUGi8cJ3YHxmLcfT9JztL6KSKKjCOILgRRnrKzXbm1Bvhe
jLx6+i75BTktVv9Q8/8IrpQcJAzf5zS9Pxd1uJLbQ1VwPwmHAa0bAOycwn1C/93d+pV02kxcXYdI
aFqHVePjVS636j5VCl/L9FUzR6yK4GVzDyq1+jNn+5EwAkapred4MCd028iGyPoEa9SW+rg6ss4n
PMGe7SyZJSc2qZuCT+PkxWZgoaMl1O28hLnqxKNyyLgmG/NIr/dTmDUSSuX0WAXf6wJUz2q9AqnQ
PMdHSoQMYriTZ1sPtiqDF9P9Q+ylvhxzBvM+DZYmqFXQf38eeGY/k3/4oTdGRB/WNERLK6U8aAu3
Gz5JS94yL8B3wU4CdB9l+KRYk1iOrBWAljXOj0iFdn9oDsW0HjbUV47K/WaUUVQdd+FcmW/wx6Ot
1/sXI5LbuKcZMZqZ75dhXjSSNHOj4W2bjvbI1GpeBap5J2OVFLm9g6u3YndvzfZUPRL21COZNGe8
wZ2hPbGSMLh5ANKOB2iIt6Lfjehp707sKXtOow1SOp3bM2z47Yi/rcYBgFYrLs/iqIvQp7S4Auqe
JCbFGoiniyd2p3QQAfxQto0ANDAZaEu59ZJVzV8PYPe/hN3rzqiSYpqveJmjk+rzzYD9QmtuTbD/
yCcrpjO2oFQOLFHUtylex+vzfZ9oWANYa5johQbVu61UFoBOK4BMrVxe+lH5hS+sr36DzKHBLZqd
1bdNVZugM2BFi/1bj/aLTIstsTLCK+ut7VFPIIv0yV+Jk7SU0vSZ97JluukBRLMH7RSfYj14Uvji
2b1DRltbOV0key+T694DSZCx2xiHs71oUCtbaBOewYa4gDLX3u4qsVjFCeqTRne46KyQxqf2ydON
vSNUOTIwNF8QTegJecyH7RSsF9QYx/0sPI8Ug1+hhMIi8H3qZXdPJH0/Mvcl2+c39T50rN3Y8s/m
fCFFg+JMVL2fJ2CM6H3oHN1NXi0Yan3OVT3nKVI8oZw3IY2qWyrxfEax5mY5LfaziOPCTWqNXFvZ
XPDGwu+P6VF49b42p1TeABUN0fYY/8pLq+WoPqdpPRaL7UxLRcOXv1RVlloMeZKEYkjRFHSmuLbC
3D8pEFs21XMDqG8tzy0098NDACd/HqXPnOSJSYGTNidT0yq5Ug+E0p7rWZb8QOs1h1PqYpoZZwOJ
96gkJLyGtEhAYutjp4x3lcPpaQgfwuvzW8Ob2sQE6i6zcTThtuveq+47Xtn0/6MsjqHPZLpSKakQ
Z7ULPbM7JTSdJ6bG7gjcjlsQl/GjspU4guib5+yilllS5YcOaQJLTZfJHAuSeQqRvYq6fpKlAtdx
9fs/KveDSM1obUelALYGdCBjtcCG1liPbv0eyewRl6vfp9RTWVW/JYXyJnpIG0zU4D5CHeowNXju
tGwEPZXjKkp7vdpH0kFLK2k7gG9Ca/ZocOP9IG1M/DjkdCqKlpQ+JHDX/nhbD1Y5Quag5YdRya0+
zZzZtz/ugSzjyX5hS8/rkeyRuuYsKSzAGEKSLydzLy8PlPjspIpyp1miO5S3DXTOg9Mpv5IvJV2j
OVnWJSTUOlERnFlHIbZZizlkNUfuGzr8fZWEuyhW8XTxt4M7hb71AtOti4O6p4ofs+cbTgzwB6J9
zwqP0w03aknPYiTko2QvpCrLivpAy7Juo2a3ViDvJ++wQk73i+dSKgdEMSj6nCRfpX+ioEFPcOee
zjsIsvjY+7yBrnJHZQUNJ22dDgd9/drwveFXMSjVaA/M+zhbK/aTbPAZADm3m+IMEmcG/2KC3rvp
uViLrwYLa+qeXkXSnhl8j9Cgopxrcho5pn2m7KgCIU1UcEitpbYDOxHdYJfs6zEkSysnQu1B0AdC
Iu15E6wsK8gy/8zGBWsGjwhsh8zdTluN9FFI/mPWxNelAISJ5Tbz2LQ5q7uFpMX7Ze+rDztcSOQN
A8iZSymvljgODt2i4OuVvo3wrFCmtC8u38a3KnnnROddcgNFhxsLYjYDXYDGWPUpjgAAMrSxJ7SB
WktCI4+3R9dSOjAsRhx7rcjVMxuE4BVfFniA30DKwrtf6PaYpUDPgOxost+iqsS9RNpvH5AM5nfU
8HogTYE/OftEpF23wFPWi5RkZDC+hbx5B6GfZ/N5O5VkdviP/jP6M5QojDFlfrZRsCjfumQvzQIF
FkKN+MPBoSgcVFNR3gXsmeLDC9oWo8Oqubz6LNAZ5JzAtwoczQJLbrEO1rSmRJ3WtE1U9bigcZAi
YFkbp/B8zTO7B8TJp466P8MJBeqiUhVXasdG73n73vQZ935FBJt94/yQAI82PGSxeB3x2TYyuc0p
sxeAoYXZbqiWO4kcy1PRTUn3CRLLs6KyignGJUNMlpwZTjf7suf03ydGHY3MoXW0o0cXQ35ACl3+
A5dou8odVffwzOf6u6nyiVdg3bDDCxG3giXf/z4aP6GJeHrMGDiWAQYgpfF6tvQYMj7Th5URXRag
VbPj0Og4xCdKkJwGDf2ST/nwNombtG1nyISkAVSzaPob7lPRbczBesUrpPpihFavkg+wo3hBCvtj
vS/c8ZYBRRcmak4MEu2ThccDBpOXvcLZcw0yHtLzK26VqA8joCN0xpmyK6RVvk4794e5W63Ca49R
Y1izcANDpCiKytyrI952HpY8aIM2YmNP3JN+ZSWvHmDLuXcot+i6cHo3TK7rXLVB+vnICyJwxo6d
k+Nn0LhA9Z3bKk0PHsMC/ppnGRlHV+32rXfZpfApKk+t2wAcPAr+TxGz/oebDiqBTQ1jh1LMWw7f
wRw5HBY/OHQwYWH9T3XeNoe1g259ZCVEHhrEK4ttZc2ZWttGH6Fgv4jYHO5TkVagH7Rrz2BrlBIW
073brEKXtZfJxiY4AvMQ4WK8BuNwK2eb/oBRrzs2ci18tYVzCcCSNxkVLEBMET9DAWQ5Wkxh4dcu
s4GqpBOuepG3iPo8iknynO7zvHAhvxtWz6uv8+iMuXabwbL9RlZnGlSfWcAb+eE+zG2LRTEYkwAg
o0UtY7pV6vAu2xjOPJ3xK7PU3Rnf8ELAbabK8RIDYBEysM1TLLqKsF/UznEWUQn/NsbKQdSb7kuB
I8z8/QWzVdo+VowSNg+0Jzl39/O6ztDBrYciiWjSUTtSmJnu0NtcGkkrLq0GvJdXbOZ1WrOv0ZBY
xF+0OPI13mYl3i92uEb4Qu00JW8MuekALKnoW4rSlfr5DMaeY3LUOFz+Qe4lpVXK+BqJEn+32ZpW
4XxNSkMI9PSPxKpTDlNwOVRuTCMcEHeufjad342Sk6L8oAs7hayusGiKE70SNASRlIpHpRvmguRq
RXxuOWJc84/xTVQmFMSRJuuWxrXbUDyswsUXAYVBAN/M1srf1Vkc12v8Xxd/2oz1911a3WG+Fxve
seVhZrRpUQcHtcX8/JAX+MnzGMMjv2uVlgfXQeAMLSSJ9wSuaXr5OX3S77+tQYSUGmVxivqdG2Ef
0DDrcnwlclyceZZqPoQvP0z2S+QoSpDBiu9WhHi/mQ0roN+9ZG6xNmEDTDvO88yviSoLmRWnz8IL
nFJ9kI/IAmUrfvjJ7z5o5m9aD7Dk7g9sLw5T1SvhoRIC38MmuxqBOIkHu6rZQwGm7r26KHCCbPBi
sTJjVZjC4RHHBUMLN8RM28HHeLXqz4ztNbC6zMcVh02fAb4Rs2mV3oMAoG1U6dt8oq/R1WTFL/VX
IB2ZSeMLLd0Anghz0IMOiXw02B4D5yM2iOilkkpAnx15LbXHzfEdMudpBKuhE3lqN9V9wLTbrZS/
mNBMNLvTph2FDhCBI2WAz4K2oADBYq10ufgZDhQLPUDFgSWzygx+RzVJUUrEqxXp2qp6RvHBlqQO
xBXI+6j8F0h0NF9GklKOUutmDpyX+jFGehTKUytpfvdoBAPe7S7XKA7rBfolLP2LwzRcKTJf75zQ
PovkOktzrWRTxIBxoScsYacMGToejJRKlHvh9o1IwVBa0QR4tnQlEEovzUy2YjqNPVUNY0fHdOoP
AR5ktPZXAa0Z1Jx/0/W3bKMdFdziqDC2eCGjwJT+P7JPEP+PHi7XPCreuriuOng3U3DoNzDBnCWl
ahTOU9V/tVGViwfukfH0ejyFIeSVNjXT4uNEpXNADVNJgwmBC8K+oWiPGRLeYb4zPSZ8rVGY1ytp
415pIdqjYqRS16t5iDrrgGP4k1qoIv6MD34v5qfG7Inaaf9idp1OQtEMXne9/G7WsoF4oiyFiJB3
uPTbiZU8FDKUnBZy8T59HGSZFTKXgXQr5iRxEXe0NtF+weiw5pfMwi9MFArgcRdKERLLfqfWEUnL
t2d7kBgZeeS2CORyLP+DlyMbAFrw8vF4MZrmycrzlZDBaNbaXyocOVh4jBDf0mesi8N7b6TT9/FX
uDYNMWtL4eEqUL1FQzfdGQj81Ztcbg0gBbN935MqAByuVF0zMbZpVs1GXwgKOeVoz6y5+cGCTDGE
Bpo5WfXnJYd8F45jEtArjaHdZXAl4SFjXzIFEbe2QK8CIQ9eaAw9ASwkTETa4KScpUDh0gdma8IN
HSSQ5oOUBTruhBeGhyOskjmcBGCNb/ME0dlTNWVrHzK7FGhSx/2W/oap25mVr0Znt/lF/pCKmF6j
N27H7VXoiCeLk7GyHOSiG6ON++LUwPBBtDIj8+tIO2lngD+QWeegFZMlXJGoBOTIhXdJyh95NIma
0Al7rA94j7BBtVEYOrCcZTyMCESHg4vbrHgdQVGGBupyQRY7XqYSNLeiJvLQmvaLC/eoRW1OzrLQ
YxgQysMAUt28FPymSCBIFBpDQxmrClBEugObtQm5Qk1//tibBldYnOeytJ0gBNJUe23hdygQjR7N
HvqKh/4mqdnMEmJWMwcFRs2yVDIEdVzEPlS4xeL1Q8Tqup8qphRlOmv6QLkRr+I+Bq2uHqD8xxS8
IXkatu+dtyIrE+QpRC0feu+26us1Py5Li4DGVldhZk9YtdwvpwquC++VWYlQIQIl/o4AvDtGcKD7
EnTWe2sy9Ob0Rq6/u0rfelty6ZMua8QmA5BL8ue1vMU36BzcbkvTehG0egLatOsyjHZ9jEuM6LUy
oyJXeoWv4LT7eM2yRBaTNNqgge4TgLfRMk6ZktOADyAHO6Lq5sArVUNfkG1prr2DuVxnaZnuJZS+
Di9s/tbqMHRRYfdjXKpqkyuVvefhgVWe90brWNgLE85o6ec9StwIpiKBTHM1jGc/VyuzGhD6cPqM
P2V9syz1jHT6w4vQ8b9MeXz6QIuJFJQA1zZQiLbf4ctmg1WpMDNogEoYwn0zsU73K61L7595r7/d
4WE4H5sXBgE4G99KraTzMESqHG75LJyW0mmWEktMJCL90DCjc358RrB6EgelrKNQzKMDgovzuYZq
sEVP2yKcfqrT7wRc8dC0hay+QlXepdKfLjU5eCeelVocd+VVoA8X2gXTu6i9aOIe4c0Q1SbY2kTo
hZWe9WX/q1KkIv2eikLQ7DtDSPX7SZoq4eZX2w392buj1ajX4KhppvC5KZjEfUrqrQ3BCEQpmuRh
4HfILjX9aLXyNbQHwbIjUeF2JtIk67CzGc3Q/PwOmUpPx0SkCj9re2G8q5Hkeswm8YJLjyeTg2sw
Yix0nzSPLj/pXA2f83rmy8yMGGp+yxakcm6Vq2pvLK4WFbOdB0Zx59N/B/1NjAaRDPSi+fLEK25I
fL/NUJIT7mliaIMsChomgnHowHSR+aM/3FC7oeam6DesV3+KAu55EpOXEt7+/XI/g0EVw9RY+NNI
EuN+Wd+BEAuDdSFPMN4cv7l1bGPZbwp6WQtlhH9BVuzBmLzkGQzxQVm7iRid5I6oUYuzKGg5ZFCe
NJz1gOvt27NXt3T/b86xZKx1O6UqZ/YMLWFjFuBdufb8yZ1BfKzz7N9KRUHSY1UEp/i/dpRkmcYN
qq4/2PEDmZPAs3XZzOhZ92BAP4jFDN/UNhXI7XSb2W+6GvIUqxAa+jr9FggR57q3QdbzFuVxMeSe
LLvHfNRLoFuJXyOpwsFnPEEvw8mt2Q4EW9cFI9nyP/k9tgfzVZNPmsSQVTW7FUhPrS5EOV5oYQxc
l7nWcmAF/QdvGucm4Gt/JJIcpxKcxMuDHBZo5N5jvEtzfcwhngfGnYLt9a6HiCFFcUW32y/0bgWW
GVnOFDw5ZYPUwEy4SW7zve8n9skCR1bOmQsf3ZpR6hxQX5DDCG55GyxBoJ0V4JcFzSPRaL3IrCTu
iyIbbm6HuskhOpOLSp3zKNjfbXdYIjnme0npf8/b593BQz6wxfYAiI2W0sQpSQQB30+P7IXW4rsG
9zIwcVJLhU+zOtBPoycU2Y7Nm0rCjkZKolPvTgkUKU/Ydg3G3Lq34JXqTQyVjW+V/3FFQd6J/C/Q
Yj8jONDgPXebGN8XPAghYVJGTniqEF+meaAJ911KykS03nI6MyvOd4hKVFcRMgmvijwzCvow9Ly+
vaIX+T06/R7k504BEtpxwIdQEjO6wpzanZTiHKvq0BtsclVQS+IQYESZ1Ml/RW3CrfGBmQARFtla
odFUrkCBFkU+Kg8J4taX2QwqwnrX3UqEuXU3AN+EU8/0eA3hC21yX4akhNiF+TEuQLRHKcr/ubD/
ykY77rOU/Mwwud+gjsYBNlDBaEc0i2b5hO4VRXJLOzYwkmZkdBAwQnE4NLvz+PItRTZrDozi8WOC
PHCleWRSlTt/qiO/VXfGSzuNjBQxDzLt7y1V27UEuxO2CykMOTMf5jitBYlG8Oyo5Z1jIVmIq30x
1cPJcrHPL3UQXrTxEZe1B6e8Gk1RLQ1BIsaqTIKFLwpMTQiZaSfrSkT7ZfdMtxaVVwry6CfJxMc4
dP7xfGrYZmUEb995wpzHrBNkWx9t1WS2gFE/UXj2SrUwjXzlOBjePwy+ECQGS9SqXsj6Y3fF/GYG
9PnY88zyWHiz0VltSe98gr7AFurDfc+bxl+zHtGBXiZ447RUwx/yqlYS+wMucpsQX7bbjCXiqcnN
NPW10Qgn0UPF/VjmWCL6T6VE9e77F23K2BOBv350cwda+M0FYr6ZYIXK49PFnsTPSMt3JxN0mk53
mv0zAa7a+3qh/yBC7h6QRGbPCZ4mMbAeuPaUuDbNCok9Sa+6lI1vo2OIOZt+6+FdILrE2412ZHMv
8IwnZbS9JazD7wEzsmfulTTc+oDPnqRmFWRHYf44Lj4xzJBJmdhog4Ppqa6AnMiUZmz0D2i8asWh
uWSEYMD7HulBomWxF8lPw/2jnrOZ8cCcM+7hdkiN/JK2RcSdVghCDVqt6wQ13yMWnKQYq9A9jv1n
75uHUUVLqBRHLUE/8nnyT1JSHTPtRCcFuYulHH/VWxxnbrIq+hsopMRtG2XbdOTCxcMUkNVB3iOF
nDTrPmLI1xXfRloIX6OXh0WmJbq8yzhz4J1UHk1Xe04FKE9D+CUzWwCy3vNnvnWRvOZmXyURygou
b0BGb8hGLyf2EkoQkjW1KQ2daW7xDl75tOx9Dwgn9apwvURHciVokFT8ZiWQBsHXXpLE7OzwmzVq
cBMUQCrJc6fCaB0D5HJvBjL8UtB3i+RLZjMTNP6OilCqsmEAvxq52GcCtMJOkAXwCzm13KR3Zo4R
4RcXzOPE7OPEpjOzxqgZdETTpzRXf7o1OCHABhvxSSdHgAquUJfvl4S45arG5s5xJkGxB53jAh0T
x6fLipZrDC62cE1CWCwPCJE14Rjhb2yZsjgeLYo7TTdo7ZF+29klskFQK7j+6nncHo/dxnrAIMdJ
ZhXy4/88vI3MthufXI+wegr/kNNfHj89zJiJPA4LgYf3Y0hNz7SK1cXU47RVqsdBEpgVCvJi1/16
7LYeXJVvBg+5RJjr061Hhp6X5bKaDFMnxT3sai1rWckswmlNG+D1SqgARqP6p9lWpKQ0xYBGc0Ox
ZMpPriFu7FMpUtkWpof4+MkmIiNejLIWozoG5BDM7XWPWro6ayuN64fXzHtcgphc6KXaQ6tzMgig
+yVo7VrhbkTKKWOTdpqJfUZroBshq9ZhULkZg9WBG91XCk+9LufWNQwvctkgjlIxPMpeOoh73vFU
jUagnFDP9tOjy3LYXOVV43nE/Ol6jNVyFdD0LRvLnzR0kD+aNMCP2aFMyEdkvBKNT+uzbT6UmNe0
v2R6ZRqQhV/6pp5myDc0mGcjkXDQwyAEJUXp8HENcUW2N+Iiz/Il99Fo+vmSiwYzj42rpVLDX/IK
7cHRjHqLwnnkoQzrpDP75XmQUn7dxF/xx2F1LP8v/E6PdNMMBv0eY6FRERfkvKv7fLAoGzAvRWff
pJwaM300YzFOBJI2PFDbh9uaKPOjGZFthLHVW4Ww3sSa2AePUv2B3oVpBIaGtdvwqRuBy7ZnQqww
yEptnrjF45Vzxr/1cjJhtS1TsBjD+EIzv5g07PbCe0mPJwria9Cc00nPDvPaeEA19NhC+gLQg1+9
vzNRJRr/20smGadO3ThXwLF0Dnt/yts+oa6l9m0Xj0Kpdp/AQtu3NkEchBMlnLYar8j9O5qg11dj
JlEkOp09wMXagLCv9OuQHQU4/Jtofq4I9/uulEDiQZV9YAkHuujCVB2bknnGXXIEvdcVPR4uVch+
sVgElQvJg3nQqnNIiBO5+FSbgRlYzoLtdX/bUyrRcsfHy7tVvLcEdgmo/AoXKicsd8JGQ3CUNS4w
UG/E/AFrgK2JOQFOVtVHswi+5MAMM+Hv7GR1FL4mLLKrtSN488Jg2SWP6nknqyCMQAfDfRxv2cUh
B9FUh4Xp7hDnpnxWycOkzZOB74Y7GZCaKzJeu1eBA0YhtGfkEIXt93oaz9GDZTOVaZoF5pVuaoE/
zKEpagMqVkBNEbLhLBBAAtG+KgwFMATSdWGedze5MN+4H8FjvLSX86ODzsGFzzTvSD5EgdoqhzXB
6X2xmG0wsjYjFqacaw0xfrU2fxqdGt4Qmy/2synAGMH9oZbOr1CKUgfUMcu0OxW+4Fgf0VDNk3Ji
nKM6QEX9PK6Eo4/pSdk9gxd3Ac6j9jaWowIFt2qTA8lA9BjTuoQXdgVZzWpAR24ofccYNnzaeDpK
//xBzV1355QkrFfkXbwsCLgbLW/UOsPqVa6zFEgCMvmPXzvFmXTyOtCqXZpONeUzJgzuU0ANbEGt
b+p0vOvNoX4ztFR+GvQhBzEIZXCRLbFCKVn2M3lrMErwqSanfGvVwbHiwQWpLZByt3QQ8YsXXTcH
cS5kWS+qr0zY6qL2yXOAWgrvvb9WXM+6hn9Z7aDjHHK9fMzJT6KBBmPSVW0Qyl947fl7hWLfOxkn
tpjMF1RjOTulpnZSAJSLL2G9ArYg/wP8g4C11Mw8VnYOLME5NZbE4fNcQHi3oy+a9E53llcEeOfa
oiVQE9mNkDoDrZpnhlWoxlJdDNhbJu7KB9BwlbzU+rmif3EKNA28GjVqZIXXecHoA+uqq7z+dNNE
ledVDNQFDOQdu8yI8OiVkoQHLygMotFOM2qY72zjE8didm+hmwEMb2teKnaoC6Ddld3ta+7TpgBz
FKbCyq1j8hmrmwOD59GuWKrxycJtZFiR0cQ+gTzE6tJ+7uAqjS18yvJG/H+U/BpGwRPt4d8hpjUG
Cpqg0drWddSUliaiuKqo1O/ECTIvASoaNGNapBSWQaYIz6fvEMdl6Ne2z+Cbo+U1lAtNiwFfrA0M
/zsn5FHYWh8nQex3mMJFCzXWZiQyZ89jzvnDNH4KaunX+tBc27wc+31Rwp7/LUBSs8SB3h6rxIhr
X+UlLo1EdalCXNGSRcgkcEzWEw3mPGB6EnwiLVgl9fqoJry9vnsecjBWuIeGXPScm/+snMUZ8BxH
tTR02gZcSK0MY/FFI9fsWoPGq9gxA3bnRhSo5avRa7a3mSNIbmd28n7U5YYdXlSAZawwa77BzduC
qx3Uqmop2+fou6Lergv5vxXzrBmTjhiAg6S1Jamvdwp664Qk7YeOrBQG2I0MCMPP9GMnIrYF81Na
gMsLdfNUrua57B0D1NFhWbt/tO1o7BJJm3xM5aN16tI294ELEKOe8cyCB6SNLOg6HuK6mcWHOrEu
P+dKFVPr2r6A3e//fAdJef8OLptLoUDsLrSELwVSmLeLGW281asz/qvfHAxmQF33ccp4f9kkTg6S
IS37vOfEP8kV8xDZ9BrVLeA9Cx0aM/Zklk3ENnP8apy0GqDvR7LlpoQKFEbav8LEoQKHFSsfQZpK
mHL4iPVZDyBT/a5BG9IV728HLxCMoekFiAed4ARHo9Dr+2R/lnzW6tPwoSx3z61XbxLr73wmI6Uk
/auH0LM0UEpKfFAhP6DzlXoPIQyV0ZONZfufYUhxBSleJwHcNZWJCLXT0tAHoRL83GZyXdc4e/Th
vS9azT2JvWE4M5vPdQvWpq0Jhyftl75rqQuo+kM/NIeBO6QDWVlLFiVHeajMkTPZfyH81x124xm/
TsCbXtjx8HTPnZXqCfBstiGIpOJDGWcvHa8dzNUv7lh2OQukGlJduZ4MnU1s1zHULdLJS3LraG38
JfrP5ChWoNxzMsmViV67YWXHJEl+2a6VtqNfkmMN0pkXEcwLUuBM0atmbwHGypPGKo9I5Zi1p4Ka
2Iw++FxFY6HkXTdApDCZFKln27mMH8D9SvC+/e1sFzsIZwqcBucpvdsz067JAyiKBYM+1esvkq1s
axwH0JCXJvJj9oH5qc2sF7gq6UCNCMQhhxG/K7TZEqfFBHmnWrLJTXf7GYcNQ68gkX/iznTnn6TP
kVlM3xSNBqQQX7PX+HHcOKg8X0CQR3418RM54H7PiKIrFwIlpBXfcBRXU8h9R0PYCHHpy8pRU4py
K8ZMiXN3JKZEhQPgmUJt0+0jhMSMNVE8htE61QGA2d3Ky9XruPksqSAn0Ly6kyAoH3OBymKdnS7L
4oD8PUu8PML0HxQk6IRxgdp0fRmT4BnnySIyOokqHrlnJbzWcG+mXm7CqNN9s2yYCka0ktYjbSDQ
tgWRdazl7VN9JfrGIg9Mux4IihXXpmjSJJ2usIwPCDvFXtSU+7fXSmT2Z6pk0bg4A6snGhl0VYdp
INH77Cn66kB7CUnB8zvR7DA+nEtcUyNai3w4kMQtRlwbYuYz/21GHYX19myEaAUMKJhHjqX6BNEa
tKggwQWsj3RAAAtfYHKOT/n1Wnp9PiBpBczdvjk7emm9oJaktWqHx7vv61Ymo4LZVjRMQedNxyGj
AOiYLAM+YbcFuNwcaBxcGPo8rPocghZ890gY6g+jCfRFUPFJh0mKsaA+W8RYQQFtcPIPX6gSsFj0
eKGFzMvzCBKniT2462mGkdnYaz0VITE1Gl87N9NEbM2tZx5IjME19quS3hdLTnDlytFQlEswBoqU
F3vgMmTmdJTSZGjcC4G6t2WrRGA8+CP16ULE0GYHNlLcVCKEUJlh/6R/+K4gwCIMUtm+IzEHqn+2
hmHioB5VRjfOJ69bFigQqm0eZ2H5IMfzJ/VWpmsPHAysjQQsOrR0Su+MHgfdb2xxV7Xw9OL/wV1d
hwheejbfOHLchE5t2XptWZJKheAzUMU9XtyGYx72m0CbXjbDHunXUwzCZBHqR68A4LwFxG4Jkhl+
HB9Wnqgvzco+SavzUVdOjAjzQ/zn4Sc48igOU7Fca0xd3WqNteTy8WCyqXu+vilAUiONfiDpCBJ9
Yrde4MOvvCWVyqRP83c9CwDtmfFPT98gJLDr0m/72I7Tf/pzPAVdDzojlbxKOSCOtj54MrY+E/y6
p2sbo2KKwnYWZZczHv8jX6tc3QYb6fswXEGS8/T+YCsdjKIBD+SxN+Mec380WRYn8stzFRtuNG6k
aG6Vvxq1g9e9qVtx8yWD19KBiXeFTtjEXey+Ilm34ktZyt+ETI3fZU8oXGoXBZdld+tZyMVEShIO
YMIbHKsH+G7tJGLPZHVc0ZTUFExTtjd54yUz7L/GxxQPwzSt6A0+ZNiBOq/znCCcZc7vgfp5xfTo
GwukHW+cxhnwffB4ykIo9/zbDtWNMd++sZXq5fsdVnFlin+KYCLnAQfMy0a3xFWN8yf0WLSktf4J
Sl+zCmqNSw12PpcTfZtgT+/mqJEpjKfuc0UfukTlVQkdMIabO+z7c6V0ObX7E2V0qAK+xBmYo4sk
1P7BFGh9ErNxHmAtFVazxdaEpcrtkpCbHjPUbu3UOZdAPAgNVFA5m42gTTwywqJTSj81mY/I6omR
JRTjZYE/AbMTiaWogTQg3hPp1jqfXR7oklHv3h0GdHo8SwXmaFHGa5fx1hYt+3gkxXLzBU14dnBO
X98bsE4mXEL90WfBtA/uLOfW+TqfbLI7ALRsxsOiIq/nYqJPi9mIumh+OxcUuWPcmyTbqnkPrzT0
Af8KdK6qdS5GXEauIm4YfM5Yo6F49hfVZAxM4NQe6EX6e2gk/E58SQ2kqq7OnlQWwhIVeNWTD6LV
B+LGThMuP447i19wdZTPOTo7P/jRGqSQYoJQbu7QdfP2HnoEAVjylEOKFIDUi18G0Nb8xBUwEh2O
LUmFHqVlt4mtCm0XJDQikOtQxE7ykr9tDtceKQuBBxiP7lWUGOvq/pNGDnV76FFWMQu4c8wq0x8y
Ru07Y8wO03R7nsBNSTVUj+v1THaNWup4wO2Olo0cETAaQ3cXRg14QcvYJnqKmRXwDwz6t/EpMmY4
K5B7m2ehC3OwMI/5WcsbvgSXM5z7rLGktkKEfjDme27SkckgJE/iJ5/B0m80b2ZKCho/g//uasLl
0/lr2PGdVFgnq9kjyahPTay1Dw3NxxDoAO/FFRIUOzoxP0GbGoHJpASX8kVraKhurXPVBrMeBuPY
COR2qvDEKfSKdmCg2q41/GESCj48/nBUj1q/7WF7ndZvm7qgBHbFtQmCz68iInudN21q4naXxYqi
W49JaOBC20eFR6OXCw/zkPRuNi0vJVYJRICZtJwb48n44f4RKo0cve18Xk5uiWfH2rtS42urQW0n
3cjmLqAr9usKEt85C7dNObzNI2ykL50FWCsDbKmeLwKDfc0l8AsgqykgMlMJJoj3SBPtsFK50ew/
SSQNNsJPj2hSie3HemHVXayeVlhG0njNEwE7eNFufsH7ABHieXqIzvBeSZQd2LKixKS/CHHp5G+I
K3ITqu1yAL83kGxFW2XE2ltv7t7ePQmCpQ9HMaCTR4J2lgEmJrIfhU2clBDQqBGyEWh9ROwIVDm6
cmsLMNieytftFM0v1F2KB5m65zmFB6vWY7SlLLZfwtN51ArnlLA6PXdubtc+yrV6psdah6fgfHjg
Q/LLlRMqPTRts0g1SrJV+nMnt4bQ4bZCrJLQGHGe1OrzAFMR7ynL752tJXBO24D5naAT3OWk/BaL
nlNE1ukyo9b0rPLgTwWUJaitMXV5a54oL3HOjuC26fwMiroCvNrBAVwoaaeIrh9arNCexepvRUBN
VPWcxO0M7JB/81EXiID2IgkfZKl52nFGD9+sZkooVYlMiv58rCHTD+7ISGC/uFRPxo1B1sWbqgIX
mtONndi6idGl2vdr9CH+xGjLtkosJafUj9fX5mS6lJiu4U6FGJw+t6byYTDdzord2h5AQ+NqPMLN
LLBV5Xyy3eLz2LmX1jJJqyUQU+7qDdFk53LLKno9eiVGOJWAc1OtgkPjyrBKFW6uKHAhtKgTcKhK
Ke82SGngyzxL6TbpnPNnmKiPWO4iJPxWTDbGP+QWHTIjhK49kSaQVrf3rAFKcMr4zaLNWO2ACdIX
EfqkxOPRxNS56lojF5lPyhJVpts7YSHcLSdeBUHuE3KNMJeMSL9Bx4ramAGAxEwnq9DnfvOmavDb
XBjwAd7kY0/X68p/CXYhH6kg/FWNJakLMEVTv/IJWyYg8O35HhJpJKIJXV8KOV0QkSrl7SQogcGP
fL6uIxSIa2nT0Tl/W6oWkOsGJ+twlKSh6LECPNOtuZYeFQGoSFv+v2+tQf71LdIVaA5JD1ZswDRH
Sd/LCW8/uQHwLcqZsDshUOq+TDgw5MWfYIRto7cFdva3CbEbHSSOAT76wwGhb+4lYJKLftmKZMsj
2J8p+ZisAnTsZqTsBFe7rol/UAu5L2InotMjtaRerLbCJS8I+/6FpFOLsmDxKYmyzhzSqcZym/xn
ulgy4Ecp2/WjZef9Jcc6TM2vqrUpzG1itOwL8ntpNPdpq+Yu6oSaQYJyNOv+GdKDeedSHTeFsF3g
sRdfl523GWmo104f3nUzGNCl/TUiEECkBF7U1A3RLrRZv9rF9bKMZwfj91IpSRO4wC2B56SkpRMX
OrPB9LJdKZJgQoD9r+h1nJ6fkRxU6x/2Sl4HYcDGUeHTrxKRnoAKOcSys1N+SFZOGXCUYPean8jL
vqhxm6EuLCilJ/plrvoNnE1ZARUL6I9kR2656uxNN+W+tgLTCvp8FXfx8S0weem1ftKtqLICstXA
L9o2w3T4xZ50+KmNdbpG5pQffTQgf0mQmpLcuEwmdpOa4O5ozxJpP9v69TsW7cfQaVFsmSbehZcT
EO06WWbrPUhKvTNr5QnLqWSWsQlCtZaahGOwsyqGvW8+10v4ldmmKgfNT5uFO5DFkYBTzk48wZpQ
l3EIbQzwwZ7UercfoscD29G1rDOxWSE291UbhAZpIbIFD6D8PQj64SLudpq5e80oeLghJ730wGEd
11Q/exwdoaV5l8O0Zu4pArn3CUxDG/dmITlpJHKpn7RTdvHhKdlKzD+Xwdt0eqiBqr+168aTo96a
xfnTreoZCucmCRgwiE1vN5lBURfcUp7QpBQIWW6AOXuHqf47a43m/avKu53Ix5KJV6HJHLZsEemS
oQZ0fxoyxGtpxdC3jf5PPLl+rDa98zk4TCzAqdOx0LRyc14ZXnTrX9oUVF8WF22YlE1ilVC1jM40
isCXfRSeQJB5pm6/CU++AXAsrQZrFOc9vibPqvF7+Ccaw7s2GkWXnFAprbwEHRgnAhyOdb5nu6kr
jPQKV55gBWTnIg9oUitHqu7zrw+SCCJqrIsp2H1MStDu2IvZ59SgJdiboeStXlHBamTIvtkc+bUk
s/JVA5xDN9XTWgYgVxcGZdojr2nEx510VSmBT/2k4RL7+1XcaZnMtGPzMur8930C5FPVGIW3hxH3
zKFx598UvQKIZnBbfz/47Lugl1wZoSG8H2jfn6vReosDSkyfY2L9bxY8UdzzHnP8imYqSTtzcZk4
5pguIJDF9g+RUtPZdl4HH8ziC2Xu2DH+z6Vnpov6QSe4DB8nS2tVO8WVpst6QHyP5LVl70IyqLxT
5OGNW9Usyi8ZShudYScd0htaraKdez7QMX+levL7Xv4dETASOTueTdtD0pR2f4ow2R1wr2H5/qmk
45IRMZTLTMqDipOrcoFQlJ/mIi0Pxv5Z3gY+Gkd33meRZ6OQPdPOhyw38RPP1lT0QkLbjvcwAuoE
9a9Td/W0brKV7Dh9P6ZjOxbty3AL8YOFxTWHX1RkyxdOq5GGKfn1RE4HT01rOccjPJl4TAeTFapD
IxXgRw8nihdEuLw5SPNFG9NCwZ+fdKNYB1WmzUEzZ/nJ+VlCGFn2XgO9lcz3iL+QOsxIh8sIe+6i
+2zARwnxo9siy07ElTQfY38JZFXxkGFvmSSV6FCz5VSkaMAObn1LsJqgP/uiVkrESm2tRxcEKG8Y
UmXDKSyumJcWHSLzdruqbu2RrAJs1bSARjp3vpecGdb6fgDSZoISELtbse1wMnoMnfKj46VSqtKk
frDVk3cdLq7yc8y+7xPZQbRTM23JrqXUCW4QCbFHPOUuq6gcZoyfEmrr5Zoj6UFxX2deLCFcFDts
3oNk1K7b/SdSD2W5HDZZ5H8VCP4utWZ8NA8sVyBkI1X9ChqI6/FI/Z3E2vTNeb9p/1mB5kAERgzV
YpTYmNTC669HlbJpgaoirGWvptNIqQJq7nHUuMvPCwOhTbGSC6TXZ7nkJrck+b1lGX+qIZag0h90
2l/hRwUvueTpyWmLNVWN9asLAcR6tvktqKolvWnKnAmi8rssa8dJ8uGcIGeehpoSNcyHSLBNPBna
plxbL9r1pgGVZ4YYPsoAUYwXTrkBme6feyqUP+vtDcJ1pidbhdbv5jjqwJtAOnVAD3CTJNsaHVP9
hRCUmZXsmXQYyx9V6Toswze2YakYBpExYWnE+1HrDyAZAJiJ7Su6kerJobiV7gEyGOn6FVGXqBZz
Cgbb1IobVie61kKXQXalAgJzMOZssWW754mECyAyVg6YjZGLJ/0tHpgL/goczWVUmLycT60jlBTX
3e007yTXzK1tcZBFNsLGOzWSPUvaxXzpgHUVA7mcfshkLE7rYSScR7nB+FkjuXoPSjDnmIMhvvug
mh3aAdI2BlBerQgJI5Nxj16S5jwX/4yX/qsz5Tgjf7EcuAc2b3deHXwIqniD47zis+90U/kSwa7L
uxSXGl10Zelwu5Ua1kPezBg/EH0eWQKWkpqb4XnZmnTKSVRzgKprkC2SabLxznTgakNHbMjU7g0O
xU+RcgIz2Cxwgcz66DmIUOTv6k+QffmT9AOcRsTO6kp1oSeLHKCTneMcBj8OtQUYb09O2pZk4KUy
3f7WKNVefd3231F87F7E55KPIh47NPl4hYWUspWK/ZTOBcbRlhxXxI0EToq+PkMRRjjFIwnn3zre
/4Lq7avS6Q37BamuQaXMx26icxHwjqCQu8Mll/TucQeRa3YLo+RpMVBrREkwBiWt29YFwu4yNM7k
UlqEjKI5PK/KdtVao130wtLNmZ88daiGXKgDcunyaluWmbDkH5o6nKcsikkEStX08rdV7Pw0/EnX
ZbJGnnxaDP3WxyJD89NUOcH9dIfeBcwccYdVgpqJeCC5ft4Gz+NvoIu64nixxYz6IZRXtaTjnVGC
lAcm7kzW9PMYb2GJmOOiQ+PVt8bG4Lyqkr+Vqm7kM/hWVIoutmeGXUw4zlrHSXSfWl2OdwC1mcCe
8OsoP+ZysN/3aQTnsaJ+jsfNscnmMvj44q7mP9VduLFlGl6pGfKfWAH6PReJyRzsTaxY/Oar6YbU
7qSV5eqb7mdd6bzRurBlTJEocXE4SCkFIykffouJeMvWhLg7FAA59YCUVi0IsLewtEmyApEoz6nY
QFL8BeSqa+bvdyug2yBT2lt9//13mIiBE7M6/msVGqtctpaUcedYgGIjr3VV6oJ6G+dpcguLzgs3
m5ybGhNtfgRPngLXssch7oK8M/WSnahLKK7/yaBm2RJgfuNsqFNQogRtU6zlMxWnZXXGXsKXKT4F
esN7yXkuYf70oQtHtOUWPPjnvkKJkgkn0ATzYM9nq8WlrR43eK7pM018A5JkqXKXS/dEjyWrSN/1
RrlRjREQv2JKGqJmC4abBQpnscIrHu4Fnb8LYFKX57bld948zHo06ShTU9/Pa5wLdDjdMi01JJnp
T0LDLr8fHnUnkhCOi2kYUxUGQEJ+I+wvm4WpzhQGBoBGncpeisC8FW2uzQYTU2XpvrA69J42v51t
X9QJU5HXDb9OUPU5N92DhKVPo9YAVvl4w63nmwSXtTgaUjMTFZw17lGDTRCB+9ILg0RYYmS8Evil
XepUXd8tQknfQf6o1tl2hzi9qvk8GepwepuqfS/QKCnbacgm3XUQXMTUwhTBH8gZz6JD4hIXSlYG
TmfZ26kR8zKXCm0VShLQQlkyZygsxMD36jr3p69Z91RhDYNLBy/rnq+msB7xel6fIlqH+2PUXCWi
izp6fQXCd6hLcO+oLAbD9ehAfdIYLieYOKWxwUMHpGMOEMwa6JEuIczW/FlEvmTjiJ0t3DgFVK0P
bQN6+6CLVseuvOghKp62jRPkxEWJUurri19zal2Qu3JahKrKhgkvjoKIrktXpSkJk4LlntVHeCLo
k3j+KV2hYXVU7AgHF8nU4dDkhHFgcw20iudw+NOgfKs4/kp/55+V5zApTm2famKbBsSKQqOjZICe
en/MVoBDYA4DkfF6uQteaO/LM/xIpuAKvIeCgQ+6aEnz3b+rsqJXdfRGzHHml0e0BInLs6J5G11k
neaAth/MgQ7aSU4otbnJVNvFeAUKKz1y6QBJQGS078sByZOTth28ELze9RvrRI5JVv/J2R1v0s6r
Z7lI6j6to/DegHARLO2EhxpJJG/7dC12OQs5S7EkO2OS8bk62AycmtmdQExcrw52Zvlq57fc/r9v
+3Q2sR0ytTF5t/CR8VE4N+Q+N53WDVeafvtutwT25YkpWNuOYeyFnYUeMOsGc6AXfw3HJjvrkjhE
tzx/nmo+sJzcA8W6CMFc0Nb8fXtenKUZ3wyZ1VPy4vynebmHF4YDhFVCk5uBfjkNemDEyJ3pw4ec
6DXe5nku6Q3LD/uaTfcL9WMNBhmCRmF9B85VwqDYgC8Cgu8rvW+3eXV7+zHkrIMBjl2gHu81lAD1
rK4u6FaBdv+TKRWiTiorF05xfNKWtCiIPE8VUwR1YqM6Ze7450MyLykbJMM+T2SdDUhWNLrYylI4
UpZ7KP1RI2KYo+FPJ7HCGKk+Ch7IG2VypAJkELW5c0VVlh0pnCj5F6cqVEKSukE24q2OoRvGXQz2
2D3BqGhLhaXzAIBCKKfipSJzemmmcFrlhRnsjZrNHIBavnrfYldGZDpGmczaVWAPXicyTM+3wKV9
Xf91doRBy3YQYEeCuxOzGpQOjc6Seh4+nk4/T/fOZWxUa5LBdzu8rRiWjcSGI5fVXlGQHuFwir1p
VUP5AOfQzjVa1ghOM+oLL/9XUGAex6o1fU/JUeKXtcjghHhqaAu2orn4GAY5jyJyGU1OCGugMMcm
1kxpdE1nuu/uv9c/m8ERDlvaHfzKi8IKYUClYLNlLhiNuED0XKoqCFFs24da4f8B3vxEhRrRQkDy
kVjMSAg3VJPKP8jDDkn57GLnP38BgClBUq8u6EX44ij29P31pjFdkdabiYY+8vYgUmJEaB1txCxw
x5pj7cOv2mZPqJH/YDqd7VC9kZm84tELFtHf5Qvdx1t7YFXuD1V1FM6zW5bz1vssXWHRi3gq2jMn
iAEO4u4W+32DiIX+fWv/6PN6CUfcFmMfWTeiZ9q72B/xGsESyt930WHUK/tDsg9iOYNUVCcSR4PH
6L23209g82wQQAnTdb1ZJL8q62/x4u0NqXZP8CL36kO4Xb/yShqOyUQ1MYp5NEiZK2y0pGKLHPTj
z16UGiekvdNshTnH3O7vnqyeJrxGJu23rdx4G+yYN/2+gOCyPuQE6ps0PnmqXfsxpwO3YdWs5PEW
gk2/yKmUOxiNPIblZWmiMt/JxxUq6vO/KzBFxDA3v7qP+gpAScb+6mhVGiznKaUWw/Obk9qlTbVb
nIO+enLhnDuYcI9GD4Tb4wNrbCr8BHgsoRfni1KR040V1j++4tJqbZQ0BDUOzHeciWwqtCTlo0Sm
RB6yTUcNyJXmqLohVbCBk36X+IaK7wt+/1XjwJfsdTgRXehE6ZNLGoE6Zs4SONVV8D4MjuplkD8+
Q19d3M3TJ7DzBOyHJKomBPx4AGLPnHA58l6+UDP40lzZbLdrn1Kw+AKVLgafT1i6Xkx+Y2BVE/jp
jxlYzjX1CSP1mq/zrekswBfmx/by94lCseDSV3ZqbCJgTMDUVou8XZ53yzw7kbNtE3iPO0BgS3KH
sY9OqNhpqGQ4Br/Ik1Vl9iBMXVAyLhfot7e4gub5blF9gQTIy8r9F+bbb+WTApPdCdoVCU2FPYa1
EhAfG+H3U/lMLviTf9KYoOF4jmjMIc6kacDTm69Nxj+f0vsccPh030zb+CxRLto0rABXokgbjoQo
mc1/kD9cH5fBs30ecjmaTjE7j0Sob08N0aBCuM1IxekB9zR1IoBzLanC8gxHTyRhA9Kjzye3/mCY
DgRFsVl0Yxr7rg0W5f1QHhSJe1D+b4RNSdELjAsJvCnYRjh9R4JXJmKiD6yBF2anT+rST+7mcWAR
XKNP4UvGYVnLbG9iWR9OQlrtPDjwJWEwR3u4K9xcXyAFdLfrbe/Udm8npKfE7rzlOVcNgcKkDVfV
2LW8agNkbXwQvr1XM1xGV6eRugEJPGjjBiYNS54cb3xgpfDL3SXYYcf9vzLXlrUDsqt2JVbOMU4+
YKfvqnWqpy7eHsRu0gZ7DZf+5f9GO/OEyqP7FgZtDRcxgTBwEpp9dyDupbRIRSs6Wcgm8nxNrtnl
yUySh6CWiGoLHRBF2BdaEHrwGkVHQAmcbb+LNIf4RSJ1rn+6mopka0rdnWhiN9smd5AoJ4lqLh2j
ik6U4+yhJxoLgT2kSNwPj1TdnO62PJJ08o0XL4HyHMxWOAnt4iH4zHazFlAqQTCecYh693d8aQjc
Wwub+pQ/g3AOgzmwQDzXfMwklarzBY06IGKZ8obwJauhElo3PlWn8ugWQPH9TrPc+Doh2WBzmvX6
uBRoTB4rchGAYBf8tCcKgK6DLOTr26buoEf2A8iQ6oc8WdFBYXfDPsw8xRSg+wcXrLeMn8bfrJOo
vbEWBeg6E8c262h9FgmmKipglPTxOBp6a9KTNUlsaa92Djml7CITRkEN+a6o8JbHuk/u98tVQgcw
2paXtyxhyAulSi/bms8rBVAmzgTvh8pPplCiNMQcpl1jX/32KGgITXxrFeqDn0FGIwGjV7pI6osO
z2EcmUofZ4ZCKfqta1fs7Y0yhJypNJf5NtuwZRZrPGSvLn7StEtPHCPA+UhXc/etm/1lDQUK2kFW
s+HWLmVbXU03jWQlah4+3LbeerMlhz2pb2ULjSL/thlfB4vbnBb3veBa+3YezvihRtBk0xOyuL8d
Dj81pLQMhRXvRijpEyN1wZQQwe7fCs9/d+VxIbtDcQ4vujt0jWUkF2vMDPdv2x+43CUFSWQdASzm
4WZ9A1Jcr2c/nbhpqTqw1YDURim8kbvu3UYyAJ+ol4Yct6SgccRAKn8OYIqdBf2Ns5k/X/dx+JKF
ZnnS+n726uVQ3dVO8hJ6CqHmgkccuCG3WExksyWV/DgdOqnznvdzl282Nz28hetpF4OnoicOu5Ip
7fAAgsWqdB+S83WRrokA/+3bXzSThXihmhVzWRXw2Eok5z1r6oCo8WYX3WFZc5MyVFNTgko5WfR+
MEF6e+CDfGVfYfTFvQEN2aaDkrNBwcbPVQOdWQWJ6g6/07axFxSjsM9dSiLqR8BDM0bN7FwKY5io
Iw95fs4gPff3voSDKyDR9TWMSCARVw1Bx9gXJFhsVuPcZgpE5hye69e2zcpMV+aTyO4EI2/uBPN5
SyUqBlQsnvX7m8bhY4QsFWhni2HHmwvEjtRPz0uWeGJxOXSi0uOTMDRbCKhSUafPe/QgGorNzleI
FGJfd4HrjVv/NaSL3mlvehthXSdc7ij6rfPdsfZGAWlxdfna1kWkp9UeHqwnJRb/v45BaGbUIWaH
i1XxrRxPfY/NcGPkVY5jNRIviLxoNCzdi81wChqlNEbMiOpNX590cGUXV9MbHHyBk1ZYPzlf5c1N
jfNtr3vpOOKzFYDPwUeyXoqVvlweTw81J0v7gxBS0fvmcqhKETb3jIwNyduCBkxed1CKeofqSZ6M
HQmG08hm4I8dZ20LeWvGMjLnxPps80ejM7sq6qC43epV0eUCFOuFvarWqhrUrJBjRc2x8zDk/PHs
IljHt+CFIDgDGzkjoIRaf8SnQpUXcc+VewIjnSKz4Kp11STQn0c+pyX2Km8T8bb3BFiqC1l2tBQj
d4weDMkkwSzY9t9WcTvaOdQwDwZ7sOpSVLiJGrSir/AtUyq7NIf8krQXmARrWn4Vw/9MHcZkvgTv
qVbA0T/fghf7MTb+5YzAo99NuxEKa42rlQvsMtpBeQfB62OpWLmGZfspBm1KYDfsykQI0VcTxJUl
/MCSVAqgco9pblwCFbGCzTlZ5N2JO1VoEeHxmybpnarIzWixLewjhl9x/mmI6NsGzp3m18YP2as2
I9ItcP2SmLJzw8owKtLixQDlKGV1BG22BrN8Ta535rTyvx8Kl019MuTRneFXi3vPUTC2AUXs+UiM
Ixt2yKTExUEidoB3mcAkrXid3wkbuDi/HYwL7ZOhhBf6rXRSPhnTbZhbCBtQr3NGi+PtS+BnwczR
nCpoaK1DxmkyDE5Kyp8ZkqpRZQFhc8kzsEEKqFH1kEYCogE4S/3SvSmAihfUhoDRDOcALobipXrR
EH42kPtxA/g9FWkWhq8aZVvFW2w0DKwnQhSrfID6ATO9OOKqapbhjz60XeCSWpdO0maMCOYyrErm
aGQSDcdWDJt9oQUVTTZRkvRb0EhQUmMFNfSAIs/rdxI/bMwS91lPxRjRSUUBjd42m8HwVQCgXJnO
XcJutOhwO4wFapdw9HkM6xFHuaxsJOp1MP6Dubt7OWm4SAC1Fo9XIB3us9YVa2Z+GQnhyv32pyys
QrGT/MAfrG9OW1Xdd4h+NDbsXczXceqK4OF+jAdG9uImD9CztrtC3eIIAGP+au02cvmz/sBl8B65
YPqqbfimpKrUT/+MTHcM439ewORV8wnH9EenR1jxdJUfqfxnbYLjURr7Z+2t7+ckBy0naHG/fzr2
FzzBbYRt81m2cpXcBMemL/2ISJXgQfkebnoBtxwqJmeNWny8he4WkbXa/kjrxiLZDQOTMUIYA65I
ginx7DANvi0L+pS9okqLrfJpBgAr4/bejUO/UYrOBhKW/eqDyWdyxgbc/nnX6DvFhqguU4iMsSlq
FF26KjsOlGosonMdnaysofVynEfu5Ed7rDxclWYm24qJtQJhcaSTmpFJS8R/owl7T+Qee623mfsH
3FaRue/uxn9ozZxl78SFWPgqtBxqWz2o1ID3+Ev67OGu/JJdeOd3KnhC7F7XyswMtkwOAXMPFxtr
Lad97oQq7xTsFjFEvnykT/vMh81mRMojUzr2k3F9NfzT73/PaMMnz6dVSulSabXKM1zSCKfqHXGv
3O8dEYZGzPg6aHrLkuhsl7zne6qyZpnFZdTzgAXWbuQi/2v5GSQIXSzzHPzybt2g+WspKZNcp1av
9n6Dh0LN4/IdVHr5f2oZ7u6I69ERlTVVAJdY/K3VnFeoxaaLFywE0BnQ7PuIs677q1O8HGK/Ki0y
NHuYV211zGUIrWjXzpw1pxKNgouwdKCHgLicYIFG3yKKX3Hp3JLLNSjEidjWucHqj3M2P701O3cG
CQV9p2nh1+RdVUZMWwt4387gkANseTRZ9Fn5b6ojUUO2l9Qy81exi9qvav1Tqo1AxNi7o4L4snGn
TXpqwVsIth/rtuG/h+LzMuI3/QtSjWLQsDGNqn9oJXE0wEMuDKKYCubiQEovvGdVY+6FPiwu3H5N
JV3kWUFkh7P9c92YtKVPVts/61Qcj0wlyBflLK81+Va8BVPlM+uQD2B3uV5jby+M7TBWYeZaF9HD
WXya3BHTEv7aELjlEGK2242h+3zhlbc6Ee/K67x6VaRvJe3MRYh7x3TwCyB5JNugYdmtUKKjq/Kc
UPvqZmY/wsxg0l96nXA3VCgBD1h1jPr6xL67kfCqgbyNFkDJHDOXyTghmfJO3C3VIQdrHhLOWQFU
l4GHtKCWMAk5pbrH+sFmKoYQnjPXjtyBxpGuWYNYKHKJs6Qhwr20puI+nsuSFB9xWHcH2H1u2vFo
lxkW47u8voeffXVa3hUz+IPlMZoErI0xZ+ALu4LGRFuh6xT9SY/P/hy3dnsXTugOscRqZ8diDf7G
BVq0xVJuPGtGb/C/Bsa8vht5q5SqnuRdl+y1hD1nK5K6ZbCqiZL/Y3LRXl8XfiamZvdNJDQ9Y/8D
lGJSp31X7n5XCtbbS5EjX3Gjzft0Oe+N1iz5vb8D/OwcZrp2XZPANRmMGVU+l2uhCxsQYA8fW6jl
JOEZaHsenXWzq2DLE0MUiAPaV8LBgmgl53GqkXquv4nD32oNaVRs0KIny+trXRd9dXp2OA4LrB6j
PNgwThaxm6Tke6T7waIStSwmGTF/cbveOIi8QqWpjGZVPVFHzJMKqa13CiH3t5jsTUdMCXPh5TQX
iSpJ8RfQ3o363/ijHW/B9hD1xgKOhlkXmmz5KDcbIcfW0TDTbhXQ9AwNmXkt9ir1Z16LbWSPqQGw
2C1+9CBmxmug0Satdyo4T46Pr76gbpovOC3FdqGERkSM0M7tgzfGWOTYEPjSAKZZmwjCO2ZJv/oA
DFKr5Lv8x1pTDpAdibiUdeJQL7qJwqB08zTqQ+pNUakENRM+8jHk3qK+n7Xt2Msr8tSdupcpAz3S
io3T/00g7VLNUpXcBSK3PkXu0gGew/lLViGD9i1L0BGfOvOSn/Km1KeBHYcz1ZybI/bIA0AK6eYe
t8/p9pCw1onmoKZO1N9cIuo3BwxJNkcvt1QAsHahLjFNssQGb4rnUOc8NNBsY1ZABfQCq5nrV3sT
JYPB29eYWeji6cyctzUEIaQ/1o9YdirXgb3qmLHcoP0jvRXpsm+/m/PZPgPm7PqIHhc3PAy1S7L1
QmYAEbl4E9NV1R0/Bq+W7mPQMoY9XefeQmvPsKWJqGViuyg5U4UyJDOnwt6/8lSBNENsne417uks
MSBrNMxKvBtxgJd4FRey5OQOwNrXqoXeQih8YNyrjCEzInbMzPfW40NmDsDpb6KiqW+VEmk1d/h8
6uLzaisnc4d0gd+mjqCodYjEGgmJlTZBBCtlkvVsixjLyXWLFXEINqH0KmoqKjyYJgnpcKGhjO3j
K6EPGaJrvk47dx/vsIexd4Vu/3m+gSWwTms+DDvwr7/f/Iep6D4+1OzF4k6czo9jIeU26OyH6VUQ
/XT9M7SHHCgVlehVs1hzxdAO2sQiFPKcEcF2iMYuCjxNX8FjqIgSOEhlWmvTklQaWQD9mYEa4+7t
XQAzAHm7ygtObd1q0OjFp1tOV4VEMk1UiVeU9vWuGj5Xum4r4+B9SocgmvgvVvHoOJIae7ndbLC0
9nEkM4mC4CKLXBeFt4mv5f0acYHlShuc3SQWr1z4Vdt4QQLDQgQzLb3GZ7Q8C3ax730S+fci6FDQ
glm1pZLDAcosMETLSrBdThtnClvXzAZMucDesBg6hWgR27dhlr/OnOqToDtb50vpzZGzSt0lE5PC
hcN35b3gR+UTGKaB5UsVm/XpoRxzpJ+iLM9lgHOtw+oNzJSE1xcBjXL1o5nIxZP6CymYc5rs/t1q
+s+3XDt1ZoX/WKrOKpo7UlxL9pnvGK4mC7GZ4w2VCtGRyhUFVI9jUVhwcQeTDtk9UVR3XMohqHP3
Jxpt8vHwk/jvvocD1PSjq4h1QUq57kx3JS2P3jrMRxMGtLbV6lYJcurq72ASF4ybJVxC72rRXB3N
ckdBWDp4O5LfViZ/iU1V1xGit5H2EiLDEkEK7/HvBC+F9sVesxH0dqCO2ZTNljlJbwFigyZriq0l
lbkJClBofAsZe3pC9MGM3onPVETyWbNBZIUa7a6w1m4pxcia+0bmVK9n0ReOZZcM7gKJlRHG3fLa
rxeZK8OlORQTMOGxPLXqP8GjYdfQlfOTCBQMJdrS8uHQ91nd175NR7GjzHNX1T97NR2doBSWp/nr
2sy7w+BxzMVf7HfAzs/DSup9gvqqlogJNZofS6nTqQH79x9tuAY1Ev6LULBO4jRZ8ENfOhlvtTeZ
PaA7hjtyeaCST8fojPsRlC5JLyhc9OCU7eyqsGPQip6F4GwLgrggmMHJrn/UgkAhCrl0GcEtaObx
BkzCm5m8hfywdb7WuxYoIwTXtAME4C4RdtiN4emj0rkXLeVR/HYpj1ihs+G34em+niMffzFQy09S
Sr+3jNGeMuO4afy4OpZukfWC7p+ew6xtx53jbpiKo2nssKU7NrvnOcXU+fsbAI22OUDphcJzMK/g
ZQ6fGZwGdqICIMFFWZ3CYejZgMmnHVY+6ssDV69XkplIaoHkmuJcRCFeDGU+O2E3bpQi6NrTH6xL
SHlH9RGvOvOv5ONJ8SroA9F5g+DosvZJK54tDJU+0PjjdMmc1JvewVNZJ3pBBGM/lv4Ol2/dLmj9
9q5Y1F2QIpLydrQf966wCOwIK1Z0EQvZ2btueBMCc2ewc480d38PIlQrJ8GVQ8xoAijnRnF87zVE
eaHto54F5v0PL8HEHZ/gfjAmbwlN13gFAMzm/zAHL0sDwsFG3+P/OkMUarToVgSnLsN01DFOXu2T
ktJXJFV7D600C2lpF0EfVQoLth2ivpV19BDHthClWsLdBGT/bM4WPxcjF7xN16jySj9pbzwQLZOx
WQ1HH+BegLXQ8sEcxXJPF7FWQSC6BLnsu+iHuTYiCB2jf3tR0Zplv9i3D/rApUN46SMW5th26o53
rYqYQDY1e3ej6GrHeknxM+kAeLHSkqtiJHSwZIl5oV/5mI2LQot6oX0iLx6jTDddgdTgje6f7cuF
naxZxO7OI0ai/zfKGB+a/z9jaezgdemUDFQH4pIhpu7B12WmvZpwPZp5xgB+w/ZFFN6zLro4075g
OTXLAprmeNLDbUGv+fj9lySMJUR5gy5u1z2wdZrFncCbq5PPSSxPygM764muf1l3R9UEV5fqBzwC
DWLbS1FCAmYQXs2i7K/ziKMRSA4RgJQx3URM4E4k3iegChkCu20DNoD1FO93HkISAQjsEascr1T8
b1ceEiveNfq1TfeUiGSvKvoQOR5fvt9sVnA5P40isdXvVXS5hF1mO7DdXbP0kpRMUSQptQMwSwDB
CXyvwCtqN1PbOyZxIT0v8/yZzXuQVgqo4otICkow6ZplcstqYCJMewuQroEeqFHxTIuZIp9pWSiQ
LBnBxaWLq5gZfyygAjoSprarDCDXLlqAAdJbMlgwOzFCiUYT3pXr2KrCJHyjTJVtJ/nUO4YrQ7+c
D5E3PXplGuKv90ZhJap12PfiWwZRZW8tq3Mv/rHzGTRi9g3VGWEyfWX1XtGyxk18A77BDTCw9odw
7Qq8cYtCMYdyO5sLeIPS9cqv/Zpv7Yej5slzifRsgj1c6CS6IkzA2PjfYMwYmbv3Z+ipQ+tqDbU/
hBHoupgCl7Uj1P6MBySDIVyd8ahAcuapp74NOm5olYwYhUftwmJx1KQ9YaXLY8PVHV8lO3auo32I
FA+KGYO9IXsl+nRqUCHMlM58DDLOjtAAJBnNSX2GX+/secIOihGnpjP6ZdUpAHxjG3W6s+Ze5333
jOWP3PermDr0NgYy/mCqqSOVyE8aCWzvnzvAAQlGWWJtgdaxEDmnFYIoaqkdJ1qLlS6GobZFEjZH
nFjxUwUSBmZY/galpclXpSasqlyJtv/9N23/AKp3UtaXJsfBiN80FO/Fgn59hooC2gElCBgFCUe5
CMohpFveJHmyXlJoK/DHBgD+S+DoWy7w7EMPwH21cMJRny79qzDzYCvF4w323EuwrI1VZ3AJLABC
0aAW84+S6P0Z+BcmxUWMqJJyI9TeEjGK+cok2UUFoZCaDHpKI7IlcugF6hpa2Zzlk7MlcwuijIah
Vyxh0HtheMaTc2Y0NcBa5V2IZaKQEOUpvg50rNqyzJ8Nb/4ZjRev9pN8hh+Yvd1orHB8Ao8jkTVB
tWw3boCx5DpROeRLAng8eYhTcLh6h+y7C/2UkREamJg2M784pbgjwkP4Axc+fs7IwlTSYQzX/qs+
ymxzNz9KzdtJ7GyEJequ6K3ecnDHVLs92x6HzSus7PnhJymN596EYzobe9+alj2zeHvCvW4UtmTc
klLwjUEmNXXUFYkK7XhAs4wRdbDbWl5AffKfy0JYAiAg0lUsdTxs4UK/1MxjpMhs1VhX+GxQsnAv
7rZkkl7BougJDlag1e63nupunAwQ+B4lOKw0zpSbKEZvpjSBeuwmKLtKihjv1fODFOtIVCI4tTdF
O7sai1P/FMKorbFHy+RcBRY9Bnh/+wHLH0RPWqkyeSg5KAas/MHWqwAvvmUZes1MoKU4Nwu69FXy
VCtlmQYAHWtGWCj+CHDn7j9b+6qLNEesDIu8KogyzH83MjmvCvZVCNr4k0M2VvNp8LAXJXUkC79U
BMzSMsQVJVVwwivaIxGB22W76Fe9feAfFjxgjzGFsLo4tVrehgnsM5GOq/wyXXUlY7pOBxUyBwwb
ZunBBetuTa1l/x3m4OhpvxVxdTweZQxZNTw+BaKIO4sFx/c+p67//PehW4AnMvrKavihYEe+XhSp
lmQSR470ziiCJ11Qq4r5e9Lzq2GVgYlpoYPWesBnsrrq761/z53rNQ0liGOWux2lf1DnEnAlfK51
tN8N6xE8d5Gtd+Zs0D+7mp7HKWjpPBWR3SqbQwu/0OWegJ8ucpBNVhXt6i4VEmrHGHZzMDoK6GLO
QQMV3yHhN5Yfp1XE8lzEIXZUJChX7SbYcNN1PZHOZarlhJDLfWCNqy98j3crLxTY9vtG9faWB7jw
A4l+QV7ckyY7/M3tOmzhU5DRfFVjVTaNpaAAq/5828SapKEgfm+aGrVs8tgykSMGslk3LkHXaVF9
Z1k6D1pZvo279BuAjr15KTviafc6fkkm7GtBXjvjXcPU2gVdqmHLGjP19+jiTW5EyIRZnis/sXrP
mmyrun5oMFW8JGkMeKQuyxPr4kKCaLVHLuYiRnfYUXo/Y0zSN8OzvpQ9YYTNKcBG31AMNdlTJOpd
/H147nfuIPQn5ZHAuCqWJBXDILV2AfSJ2mFG+EgPqRtJs4kNze7QZ1P02WcSPZdoL6n6Ayukkc66
QUvy9Ja0UKPONGv201HpxVztRQCvRNIAOjssZuE3KgFFbYGBcHOHxqFuaOg3C4yK4HRvIAnd6CNY
iU+EbDrJEE9tEU37PqHfy146WP7RsUwl6G0lg5i1suoW3sHTtNbio5pyR/hsFE+EzXz4g698qX+V
HIurxH/mp3mrkPuAssgtoUuwne6sAuDbcsaj1YY8MwI1u0YR2WPA0OvZI0E/n11kXGbvlvC/43kS
h0hXGXJLfkGJi9OusKnCNqcPMVEchd8WV24yJRuM0kfID0YyfgdnfKV0i2H5RxYPHgOHiKjrkQ4i
p812fyfYY3dWJiA13W0Pe9lWFZk+/Fk6bQRfJjITWuI1TNMmwls4GNDalmUMloTgtyZIKUWx8KRg
7RnkSfF63CNl5clLAtSpYwDvBuWV+avk/ovr9fhayyoLMpNu15IixQpMJAeey8xgAMP9l0C44Opf
k7kFW1RrMGdaPA4wDJg9r4IZFZ4fQzjs/Kk7La8jeHpjKMo+GcTcv7qnA5q5q5dK0hdchEOP28yq
/2cYACyzOqs+r1XOtZs6UCL+dvX9fi4H3jCzZ3LGSneF/albJn65icvwMBKXwrqrtAYo+7Y8WfTU
S+beuwopxDSp11azLVnpZqDMdSI97nSDrYtmpiiTsKa78mZZmOE8LcOA/XYKFl66jWPI5OkMO++B
pLSn14qin/KGPaPs4LTpF57C2ugN5MRaLrY9rhytVYM7cujKIwL/KZ29GVVzpCeX23fhyJp2Ewaw
VZV266VD2yv+i+iKn9/hMxWG74S8CTGknNeTdZwP3CrVDLcOXpCtv3UyZIi7VEaaeKQj3Ip+8fCt
sPUwruvIv5BISFT1zfpOZcLi0OYOG33OSBUU0YO7OQPLNaic67k6zLk6gkE1IegrOVB4s8tyczBt
5g7Lwy0IicBA80bUkPWfPMpnqzKlOYgFMy6SkZpPb0xN6N7gUuwzWRqzj8s0nE4965f4qeULp4aA
zPtLAMyRSUmIU8onF+mGlIkR8QxswWxlSF+6SSlr8+0IOhuX+D9eGia/PSTC7QXEJfbrjKuO0F7t
kz9hskoBpM6KRvXeoKwvqNTJQ+po725PVOu2iuFwDAGOvnBxJshKl/4tOEyDiepvKftz0SPlWXbC
Bqtz+DwwAddY4pWoL88kwNw5c0JkEK7jnJMNn5FxAQcTsy2D+gkcUL3DVQqbbYB1lXMQa7us6snX
pj6Omp8yujZ/fQ+dXFpf1ZEBLYQio7L1Y3SzA7qkEuvM5M/IFa4/DJesTrT6O+nbNkDbJQ1456jm
fLTHtq7tJA6XDizxf7VK4nB8z38wZ10LY3GlwLLCoXAzLLAY/asvKfT9f+VRgV3zV33uiaXbmi/c
88Q8UL6bcSxnpl8yRc8La6u6W3QnJeqNDyPC5QwzWa+9NV7CFhvVEugn97N+LjjrmcYJwmV6zYHx
XjbfxenpWrBbQphHwLymnAdARqGdHa7nuXDuqxyFwOFhodrME+9FRvSkRg4HtBqEbB1R3tdmmYuI
I1IOLbS7w+xBSH4+GEoz9CBPKNLl/kyl1s7T3D060zCIZIqjJkh1gdNbBQatxhxSTm7rXQF5OVKq
JhWZlQBvRH2z3xPdfeN/hB9hbmz0s+pqZjUFo9iKGKSTU6xeazSfaOasN4Gb0Fk04XN+ObAWDblg
PuekR4OdmE4ArqDa3wnIdOr7d3i+JPMfnO1ZDH7bo8mW3d6Z9Wb1HnWW5B7IbPQ4wBlsXaSK+DD7
hPxjzi+ILKJ/ZkzAlwT2mnSio4EMeIvVbcJXtzkLm1Gt/rvA13HJyL//ayDXs2EfcV7uzPTvlY6J
SPPHDJWK2klb1L4f6LkQ1zSszxccq9SVuz1Qn/3wN1YM7wUWuyfApiHHluK8x+rma35FTGVd7qQK
qWAZF8TIaMVMtdIly0TeW7q2yyBxuLb3xBmJZRmqWNfziupfklQe9L6vGAiap2uLpZnYNsl8rqtZ
VlvLGPIaKb0+/1b0VHXGi5fDUrmJBAlLlijwPbBGTHGKfuWNmXujdblVfmfI6p24svK4x298NKM7
GG1gVgeHKbmfw+XMolu7EH10/MRUF0DftCkillIzPcJx168gjOghcpC3WWZgNEZfGsyfK1aUlsTU
TQHjWumL4GcFUPK8CJouNy8GD1VaoUPOLphCkKazrq0zC6gAfI2uNG521UBbh4gPlHTSdFPoPGVg
gRw+xs4PONEqnTKhaMrSIB809BdISZhdR+MzVVuE6Z9v/ztfIMoTO9nRM0waCQGO/ACB0De4TJfA
YHgb6HcZiBjVbKnFx7GEVkltv5d8XVQm2w==
`protect end_protected
